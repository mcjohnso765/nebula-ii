* NGSPICE file created from team_01_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

.subckt team_01_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113]
+ la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118]
+ la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123]
+ la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
+ la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68]
+ la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73]
+ la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79]
+ la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8]
+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95]
+ la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0]
+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100]
+ la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107]
+ la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113]
+ la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11]
+ la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126]
+ la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36]
+ la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42]
+ la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49]
+ la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
+ la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74]
+ la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80]
+ la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87]
+ la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93]
+ la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9]
+ vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XANTENNA__09523__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09671_ net987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[22\] net945 vssd1
+ vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__and3_1
XANTENNA__11834__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10764__S1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[11\] net663 net660 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13607__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08709__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[19\] net662 _04890_
+ _04891_ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09531__C net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08428__B net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08484_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[23\] net886
+ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14017__D1 _04152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12830__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10841__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12665__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1071_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout427_A _07965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1169_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13350__A team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_134_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11397__A2 _07696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09105_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[13\] net665 _05425_
+ _05434_ _05436_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_33_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1336_A net1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09036_ _05264_ _05265_ _05302_ _05375_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11301__C _05154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout796_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold340 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 net1956
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold351 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[127\] vssd1 vssd1 vccd1 vccd1
+ net1967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[30\] vssd1 vssd1 vccd1 vccd1
+ net1978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold373 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 team_01_WB.instance_to_wrap.cpu.f0.num\[3\] vssd1 vssd1 vccd1 vccd1 net2000
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A _04648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout820 _04632_ vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__clkbuf_8
Xfanout831 team_01_WB.instance_to_wrap.cpu.RU0.next_ihit vssd1 vssd1 vccd1 vccd1 net831
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__10109__B1 _04678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ _06267_ _06272_ _06277_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__or3_4
XANTENNA__16867__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout842 _03734_ vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_4
Xfanout853 net869 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__clkbuf_2
Xfanout864 net865 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_4
Xfanout875 net876 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09514__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11029__B net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout886 net887 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__buf_4
X_09869_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[12\] net776 _06200_
+ _06201_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__a2111o_1
Xfanout897 net899 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_4
Xhold1040 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[30\] vssd1 vssd1 vccd1 vccd1
+ net2656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11321__A2 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 team_01_WB.instance_to_wrap.cpu.f0.state\[0\] vssd1 vssd1 vccd1 vccd1 net2667
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 team_01_WB.instance_to_wrap.a1.ADR_I\[25\] vssd1 vssd1 vccd1 vccd1 net2678
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11900_ net2369 net275 net480 vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__mux2_1
Xhold1073 _02141_ vssd1 vssd1 vccd1 vccd1 net2689 sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ _05779_ net578 net362 vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_116_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1084 team_01_WB.instance_to_wrap.cpu.K0.code\[0\] vssd1 vssd1 vccd1 vccd1 net2700
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2711 sky130_fd_sc_hd__dlygate4sd3_1
X_11831_ net2334 net215 net488 vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__mux2_1
XANTENNA__11609__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09278__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08338__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18037__1537 vssd1 vssd1 vccd1 vccd1 _18037__1537/HI net1537 sky130_fd_sc_hd__conb_1
X_14550_ net1335 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11762_ net2282 net218 net495 vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__mux2_1
XANTENNA__12821__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13501_ net186 _03959_ _03960_ net726 vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__a211o_1
XANTENNA__10832__A1 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10713_ net554 _07035_ _07052_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12575__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14481_ net1397 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16247__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11693_ _07889_ _07891_ net612 vssd1 vssd1 vccd1 vccd1 _07892_ sky130_fd_sc_hd__mux2_4
XFILLER_0_113_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16220_ clknet_leaf_62_wb_clk_i net1840 _00208_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13260__A team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13432_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\]
+ net595 vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10644_ _06982_ _06983_ net537 vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16151_ clknet_leaf_96_wb_clk_i net2661 _00139_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10596__A0 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13363_ net1794 _03833_ net826 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__mux2_1
X_10575_ _06910_ _06913_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__or2_2
XFILLER_0_23_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_125_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15102_ net1251 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__inv_2
X_12314_ net2764 net284 net433 vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16397__CLK clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16082_ clknet_leaf_102_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[4\]
+ _00070_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[4\] sky130_fd_sc_hd__dfrtp_1
X_13294_ net1063 _07710_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1
+ vccd1 _03780_ sky130_fd_sc_hd__o21ai_1
XANTENNA__17642__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17966__1466 vssd1 vssd1 vccd1 vccd1 _17966__1466/HI net1466 sky130_fd_sc_hd__conb_1
XANTENNA__11919__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15033_ net1259 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__inv_2
X_12245_ net2659 net288 net442 vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12176_ net1923 net255 net449 vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__mux2_1
XANTENNA__10899__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09753__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08520__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08961__B1 _05266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11127_ _07301_ _07452_ net541 vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__mux2_1
XANTENNA__17792__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16984_ clknet_leaf_28_wb_clk_i _02671_ _00967_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15935_ net1410 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__inv_2
X_11058_ _07381_ _07384_ _07397_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_134_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10009_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[1\] net776 _06347_ _06348_
+ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__a211o_1
X_15866_ net1347 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__inv_2
XANTENNA__10520__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08529__A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17605_ clknet_leaf_72_wb_clk_i _03292_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14817_ net1246 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__inv_2
X_15797_ net1381 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17536_ clknet_leaf_30_wb_clk_i _03223_ _01519_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14748_ net1309 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17467_ clknet_leaf_50_wb_clk_i _03154_ _01450_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12485__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14679_ net1369 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08492__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17172__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16418_ clknet_leaf_79_wb_clk_i _02172_ _00401_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17398_ clknet_leaf_141_wb_clk_i _03085_ _01381_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16349_ clknet_leaf_74_wb_clk_i net1875 _00332_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10051__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09992__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18019_ net1519 vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_hd__buf_2
XANTENNA__11829__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12879__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09744__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10034__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07984_ team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1 _04482_
+ sky130_fd_sc_hd__inv_2
X_09723_ _06052_ _06054_ _06059_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__or4_4
XFILLER_0_138_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout377_A _04969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_87_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09654_ _05983_ _05985_ _05990_ _05993_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__or4_4
XANTENNA__10511__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11474__A1_N net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09034__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08605_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] net619 _04845_ vssd1 vssd1
+ vccd1 vccd1 _04945_ sky130_fd_sc_hd__a21oi_1
X_09585_ _05921_ _05922_ _05923_ _05924_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout544_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1286_A net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11067__B2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[18\] net675 _04859_
+ _04867_ _04869_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_72_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10200__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__A1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08467_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[23\] net889 vssd1
+ vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__and3_1
XANTENNA__12395__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout809_A net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire506 _06463_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__buf_1
X_08398_ _04712_ _04737_ _04731_ _04715_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_135_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10360_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[17\] net805 net756 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__a22o_1
XANTENNA__09983__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08902__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09019_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[9\] net890 vssd1
+ vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10291_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[19\] net978 vssd1
+ vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12030_ net3111 net215 net465 vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__mux2_1
Xhold170 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[126\] vssd1 vssd1 vccd1 vccd1
+ net1786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold181 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout650 _04823_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_4
Xfanout661 net662 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_8
Xfanout672 _04797_ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__buf_8
X_13981_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[0\] _04265_ _04269_ vssd1 vssd1
+ vccd1 vccd1 _04273_ sky130_fd_sc_hd__a21o_1
Xfanout683 net684 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_6
Xfanout694 _04771_ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_8
X_15720_ net1277 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__inv_2
XANTENNA__13255__A team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_137_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12932_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[13\] net1036 vssd1 vssd1 vccd1
+ vccd1 _03698_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08349__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15651_ net1186 vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__inv_2
X_12863_ net2880 net321 net381 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__mux2_1
XANTENNA__09171__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14602_ net1330 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__inv_2
X_11814_ net2401 net285 net494 vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15582_ net1274 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12794_ net2033 net641 net608 _03624_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17321_ clknet_leaf_14_wb_clk_i _03008_ _01304_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14533_ net1405 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11745_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07934_ sky130_fd_sc_hd__xor2_1
XANTENNA__10805__B2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10818__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17252_ clknet_leaf_17_wb_clk_i _02939_ _01235_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14464_ net1178 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11676_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[16\] _07541_ net719 vssd1 vssd1
+ vccd1 vccd1 _07878_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16203_ clknet_leaf_113_wb_clk_i _01963_ _00191_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12558__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13415_ _03874_ _03875_ _03873_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08515__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10627_ net522 net503 vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__nand2_1
X_17183_ clknet_leaf_26_wb_clk_i _02870_ _01166_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14395_ net1315 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10033__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16134_ clknet_leaf_106_wb_clk_i _00008_ _00122_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09974__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09908__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13346_ team_01_WB.instance_to_wrap.cpu.f0.i\[11\] net1065 _07677_ team_01_WB.instance_to_wrap.cpu.f0.i\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10558_ _04707_ net549 net536 vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__or3_1
XFILLER_0_122_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16065_ clknet_leaf_118_wb_clk_i _01858_ _00053_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_13277_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] _03747_ vssd1 vssd1 vccd1 vccd1
+ _03766_ sky130_fd_sc_hd__nand2_1
X_10489_ _06826_ _06828_ _05839_ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15016_ net1275 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12228_ net2453 net220 net441 vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__mux2_1
XANTENNA__09726__A2 _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_121_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_20_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11595__D _07809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11533__A2 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12159_ net3196 net223 net447 vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16967_ clknet_leaf_16_wb_clk_i _02654_ _00950_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11297__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15918_ net1393 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__inv_2
X_16898_ clknet_leaf_34_wb_clk_i _02585_ _00881_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09081__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15849_ net1363 vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09789__S net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09370_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[26\] net689 net684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16562__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17688__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08321_ net989 net949 vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__and2_1
XANTENNA__13994__B1 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17519_ clknet_leaf_143_wb_clk_i _03206_ _01502_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12797__B2 _03626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[29\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[21\]
+ net1040 vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10272__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08183_ net2412 net2245 net1044 vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10024__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09965__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08722__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1034_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18036__1536 vssd1 vssd1 vccd1 vccd1 _18036__1536/HI net1536 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_4_15__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09256__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_A _07944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13774__S _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1201_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout661_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ team_01_WB.instance_to_wrap.cpu.f0.i\[31\] vssd1 vssd1 vccd1 vccd1 _04465_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout759_A _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ net1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[21\] net948
+ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09350__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11307__B _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09637_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[23\] net971
+ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout926_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965__1465 vssd1 vssd1 vccd1 vccd1 _17965__1465/HI net1465 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_84_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09568_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[25\] net964
+ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13985__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08519_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[18\] net931 vssd1
+ vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__and3_1
XANTENNA__12788__B2 _03620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ _05837_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__nand2_1
XANTENNA__13014__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11323__A team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11530_ net1868 net1157 net587 net1108 vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14056__D _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11042__B _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12853__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11461_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] _04713_ _04753_ vssd1 vssd1
+ vccd1 vccd1 _07757_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_135_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13201__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13200_ net8 net836 net629 net2326 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__o22a_1
XANTENNA__10015__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[27\] net972
+ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__and3_1
X_14180_ net1412 _04451_ _04452_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__nor3_1
X_11392_ _07697_ _07715_ _04466_ vssd1 vssd1 vccd1 vccd1 _07719_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12960__A1 _05258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16271__D net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13131_ net78 net848 net632 net2033 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10343_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[17\] net941
+ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14162__B1 _04195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ net2643 net2564 net860 vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__mux2_1
X_10274_ net1120 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[19\] net957
+ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__and3_1
XANTENNA_input55_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09166__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ net2900 net229 net468 vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__mux2_1
XANTENNA__16435__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1401 net1404 vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17870_ clknet_leaf_95_wb_clk_i _03545_ _01810_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1412 net1413 vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16821_ clknet_leaf_125_wb_clk_i _02508_ _00804_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout480 _07949_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_122_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout491 _07944_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_6
XANTENNA__11279__A1 _07042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16752_ clknet_leaf_126_wb_clk_i _02439_ _00735_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13964_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ _04220_ _04228_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__and4_4
XTAP_TAPCELL_ROW_31_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15703_ net1200 vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__inv_2
XANTENNA__08144__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12915_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[18\] net1030 vssd1 vssd1 vccd1
+ vccd1 _03686_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16683_ clknet_leaf_0_wb_clk_i _02370_ _00666_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13895_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[2\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__a31o_1
XANTENNA__08695__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11932__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15634_ net1234 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12846_ net2710 net239 net379 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12779__B2 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15565_ net1228 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__inv_2
XANTENNA__13432__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ net1027 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] vssd1 vssd1 vccd1
+ vccd1 _03613_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17304_ clknet_leaf_27_wb_clk_i _02991_ _01287_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ net1392 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11451__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11728_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] _07798_ vssd1 vssd1 vccd1
+ vccd1 _07920_ sky130_fd_sc_hd__or2_1
X_15496_ net1289 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17235_ clknet_leaf_135_wb_clk_i _02922_ _01218_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14447_ net1382 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11659_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _07813_ vssd1 vssd1
+ vccd1 vccd1 _07865_ sky130_fd_sc_hd__or2_1
XANTENNA__10006__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09638__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17166_ clknet_leaf_6_wb_clk_i _02853_ _01149_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14378_ net1349 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold906 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold917 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16117_ clknet_leaf_100_wb_clk_i _01892_ _00105_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold928 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ net565 _07704_ _07733_ net829 vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold939 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17097_ clknet_leaf_10_wb_clk_i _02784_ _01080_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14153__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16048_ clknet_leaf_87_wb_clk_i _01841_ _00036_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11506__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08870_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[3\] net650 _05193_ _05197_
+ _05207_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__a2111o_1
XANTENNA__17360__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1606 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3222 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09580__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1617 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1628 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3244 sky130_fd_sc_hd__dlygate4sd3_1
X_17999_ net1499 vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_105_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1639 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3255 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12003__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11842__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[28\] net687 net670 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__a22o_1
XANTENNA__11690__A1 _07553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09353_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[25\] net673 net659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[25\]
+ _05683_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout242_A _07870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08436__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08304_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[30\] net966 vssd1
+ vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__and3_1
XANTENNA__10245__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09284_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[22\] net893 vssd1
+ vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_60_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08235_ net2668 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[38\] net1038 vssd1 vssd1
+ vccd1 vccd1 _03452_ sky130_fd_sc_hd__mux2_1
XANTENNA__12673__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14454__A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout507_A _06098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09399__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1249_A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08166_ net2425 net2419 net1052 vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__mux2_1
XANTENNA__08452__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12942__A1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12942__B2 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08097_ _04564_ _04565_ _04566_ _04567_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08610__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17703__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14144__B1 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13498__A2 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout876_A team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09283__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08999_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] net595 vssd1 vssd1 vccd1
+ vccd1 _05339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09323__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_117_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_67_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10961_ net546 _06438_ _06939_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12848__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11752__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ net3255 net239 net383 vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13680_ team_01_WB.instance_to_wrap.cpu.c0.count\[6\] _04102_ vssd1 vssd1 vccd1 vccd1
+ _04103_ sky130_fd_sc_hd__and2_1
XANTENNA__11681__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10892_ net562 _07208_ _07209_ _07230_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12631_ net2209 net203 net391 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08346__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10236__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15350_ net1200 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__inv_2
X_12562_ net2430 net212 net401 vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14301_ net1355 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__inv_2
X_11513_ net1640 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\] net877 vssd1 vssd1
+ vccd1 vccd1 _03336_ sky130_fd_sc_hd__mux2_1
XANTENNA__12583__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15281_ net1290 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12493_ net2887 net218 net407 vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17020_ clknet_leaf_32_wb_clk_i _02707_ _01003_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14232_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] vssd1 vssd1 vccd1
+ vccd1 _02255_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09929__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11444_ _07675_ net326 _07746_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__and3b_1
XFILLER_0_22_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12933__A1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14163_ net1412 _04442_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10944__A0 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17383__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11375_ _07703_ vssd1 vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__inv_2
XANTENNA__08601__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14135__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13114_ net96 net845 net631 net1790 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10326_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[18\] net966
+ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_128_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14094_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[77\] _04235_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11927__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ net2922 net2786 net866 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__mux2_1
X_17922_ net1610 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_0_24_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ _06533_ _06568_ _06596_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_33_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1220 net1227 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__buf_2
XANTENNA__08365__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09193__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1231 net1236 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17853_ clknet_leaf_74_wb_clk_i net1644 _01793_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_10188_ _04750_ _05006_ _05376_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__nand3_1
Xfanout1242 net1245 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__buf_2
XANTENNA__13427__B _04971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1253 net1269 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__clkbuf_4
Xfanout1264 net1265 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__clkbuf_4
Xfanout1275 net1277 vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__clkbuf_4
X_16804_ clknet_leaf_53_wb_clk_i _02491_ _00787_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1286 net1303 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__clkbuf_4
Xfanout1297 net1302 vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__buf_4
X_17784_ clknet_leaf_86_wb_clk_i _03460_ _01724_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_14996_ net1264 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13947_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__and2_2
X_16735_ clknet_leaf_7_wb_clk_i _02422_ _00718_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11662__S net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16666_ clknet_leaf_46_wb_clk_i _02353_ _00649_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11672__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] _03579_ _04136_ vssd1 vssd1
+ vccd1 vccd1 _00006_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15617_ net1246 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__inv_2
X_12829_ net1034 _07476_ net366 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\]
+ net1057 vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__a32o_1
X_16597_ clknet_leaf_122_wb_clk_i _02284_ _00580_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18035__1535 vssd1 vssd1 vccd1 vccd1 _18035__1535/HI net1535 sky130_fd_sc_hd__conb_1
XANTENNA__13413__A2 _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15548_ net1176 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15479_ net1196 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__inv_2
XANTENNA__12493__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08840__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08020_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid _04515_ vssd1 vssd1 vccd1 vccd1
+ _04516_ sky130_fd_sc_hd__nand2_2
X_17218_ clknet_leaf_35_wb_clk_i _02905_ _01201_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold703 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12924__A1 _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11727__A2 _07323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17149_ clknet_leaf_49_wb_clk_i _02836_ _01132_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold714 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09396__A3 _05707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10307__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold725 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 _03497_ vssd1 vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14126__B1 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold747 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09971_ _06303_ _06304_ _06309_ _06310_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__or4_2
Xhold769 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17964__1464 vssd1 vssd1 vccd1 vccd1 _17964__1464/HI net1464 sky130_fd_sc_hd__conb_1
XFILLER_0_106_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11837__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08922_ net532 net521 vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__nor2_2
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08853_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[3\] net883 vssd1
+ vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1403 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net3019 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09534__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_A _07823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1414 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[22\] vssd1 vssd1 vccd1 vccd1
+ net3030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1425 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1436 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10042__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08784_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[0\] net665 _05121_ _05122_
+ _05123_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13637__C1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1458 team_01_WB.instance_to_wrap.cpu.f0.num\[27\] vssd1 vssd1 vccd1 vccd1 net3074
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12668__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08659__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14449__A net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13652__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_A _07956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1199_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09320__A3 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08447__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17256__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09405_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[27\] net687 net686 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout624_A _04628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1366_A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10218__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09336_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[24\] net689 net683 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[24\]
+ _05662_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09267_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[20\] net697 net661 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[20\]
+ _05606_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11601__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13168__B2 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08218_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[63\] net3149 net1048 vssd1 vssd1
+ vccd1 vccd1 _03469_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09198_ net1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[17\] net887
+ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout993_A _04491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08149_ _04610_ _04611_ _04615_ _04618_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__or4bb_1
XANTENNA__08044__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11160_ net334 net338 _07383_ vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11747__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[6\] net798 net738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__a22o_1
X_11091_ _06858_ _06882_ _07412_ _07430_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_8_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[0\] net954 vssd1
+ vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__and3_1
XANTENNA__09544__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13340__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold30 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[0\] vssd1 vssd1 vccd1 vccd1
+ net1646 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09444__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold41 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[12\] vssd1 vssd1 vccd1 vccd1
+ net1657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 _03448_ vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ net1260 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__inv_2
Xhold63 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[22\] vssd1 vssd1 vccd1 vccd1
+ net1679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[16\] vssd1 vssd1 vccd1 vccd1
+ net1690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[14\] vssd1 vssd1 vccd1 vccd1
+ net1701 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ _01835_ _04173_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold96 team_01_WB.instance_to_wrap.a1.ADR_I\[16\] vssd1 vssd1 vccd1 vccd1 net1712
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12578__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14781_ net1312 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__inv_2
XANTENNA__09847__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ net2768 net191 net467 vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16520_ clknet_leaf_115_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[18\]
+ _00503_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13732_ _04507_ team_01_WB.instance_to_wrap.a1.READ_I team_01_WB.instance_to_wrap.a1.curr_state\[0\]
+ _04509_ team_01_WB.instance_to_wrap.a1.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _00009_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10944_ net341 _06526_ net340 _06562_ net551 net542 vssd1 vssd1 vccd1 vccd1 _07284_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10457__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16451_ clknet_leaf_42_wb_clk_i _02205_ _00434_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13663_ net188 _04093_ _04094_ net727 vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10875_ _07024_ _07214_ net516 vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15402_ net1279 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__inv_2
X_12614_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[6\] net298 net398 vssd1
+ vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__mux2_1
XANTENNA__10209__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16382_ clknet_leaf_69_wb_clk_i _02136_ _00365_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09075__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11214__C _07251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ net199 net195 _07810_ _07887_ net645 vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__o2111a_1
Xclkbuf_leaf_85_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_22_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15333_ net1207 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12545_ net2702 net283 net406 vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_18052_ net1552 vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__buf_2
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15264_ net1242 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12476_ net2610 net287 net413 vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__mux2_1
XANTENNA__08092__A team_01_WB.instance_to_wrap.cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16773__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17003_ clknet_leaf_0_wb_clk_i _02690_ _00986_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08523__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14215_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] vssd1 vssd1 vccd1
+ vccd1 _02272_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_5 _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08035__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11427_ _04480_ _07738_ _07699_ _07689_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_39_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15195_ net1180 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__inv_2
XANTENNA__14822__A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output86_A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14146_ _04424_ _04426_ _04428_ _04430_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__or4_1
XFILLER_0_50_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09783__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11358_ net1065 _07679_ vssd1 vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17129__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[18\] net973
+ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__and3_1
X_14077_ _04358_ _04360_ _04362_ _04364_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__or4_1
XFILLER_0_123_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11289_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] _07628_ vssd1 vssd1 vccd1
+ vccd1 _07629_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13028_ net2192 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[66\] net857 vssd1 vssd1
+ vccd1 vccd1 _02097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17905_ net1425 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
Xfanout1050 net1053 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1061 team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1 vccd1
+ net1061 sky130_fd_sc_hd__clkbuf_2
X_17836_ clknet_leaf_66_wb_clk_i net2329 _01776_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1072 net1075 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__clkbuf_2
Xfanout1083 net1086 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1094 net1095 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__buf_1
XFILLER_0_83_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17767_ clknet_leaf_63_wb_clk_i _03443_ _01707_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[37\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__12488__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ net1188 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__inv_2
XANTENNA__13634__A2 _07290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16718_ clknet_leaf_6_wb_clk_i _02405_ _00701_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_17698_ clknet_leaf_101_wb_clk_i _03382_ _01639_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16649_ clknet_leaf_9_wb_clk_i _02336_ _00632_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_98_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09066__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[14\] net936
+ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11421__A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10081__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09098__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09052_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[12\] net887
+ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08003_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1
+ _04501_ sky130_fd_sc_hd__inv_2
Xhold500 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10037__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold511 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold522 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09826__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13570__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09774__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold544 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 net2160
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold555 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 _02097_ vssd1 vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold588 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ net993 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[3\] net952 vssd1
+ vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__and3_1
Xhold599 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08905_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[2\] net883 vssd1
+ vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__and3_1
X_09885_ net993 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[5\] net968 vssd1
+ vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__and3_1
Xhold1200 _03489_ vssd1 vssd1 vccd1 vccd1 net2816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[103\] vssd1 vssd1 vccd1 vccd1
+ net2827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08836_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[1\] _04778_ _05158_ _05162_
+ _05171_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__a2111o_1
Xhold1222 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2838 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1233 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2860 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10203__C net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1255 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 _03478_ vssd1 vssd1 vccd1 vccd1 net2882 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09561__A _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1277 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[81\] vssd1 vssd1 vccd1 vccd1
+ net2893 sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[4\] net652 _05082_ _05089_
+ _05090_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12398__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1288 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1
+ net2904 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16646__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1299 _02149_ vssd1 vssd1 vccd1 vccd1 net2915 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout839_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08698_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[7\] net691 _05015_ _05023_
+ _05027_ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_71_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10660_ _06998_ _06999_ net539 vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14050__A2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09319_ _04844_ _05570_ _05620_ _05658_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__and4b_2
XFILLER_0_106_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08804__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10591_ net376 _06897_ _06899_ _06904_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__a31o_1
XANTENNA__13022__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12330_ net3072 net250 net429 vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08343__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12261_ net2452 net221 net437 vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__mux2_1
XANTENNA__12861__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14000_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] _04249_ _04259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__a22o_1
X_11212_ _07550_ _07551_ _07547_ vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__or3b_1
XANTENNA__13561__A1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09736__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12192_ net2950 net225 net443 vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10914__A3 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11143_ _07180_ _07317_ net516 vssd1 vssd1 vccd1 vccd1 _07483_ sky130_fd_sc_hd__mux2_1
XANTENNA__13258__A team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
XANTENNA__16176__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
X_18034__1534 vssd1 vssd1 vccd1 vccd1 _18034__1534/HI net1534 sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_132_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_132_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13313__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
X_15951_ net1409 vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__inv_2
XANTENNA__17421__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11074_ net372 _07223_ _05529_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__or3b_1
XFILLER_0_95_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10025_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[1\] net766 _06358_ _06364_
+ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__o22a_1
XANTENNA__15473__A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14902_ net1198 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__inv_2
X_15882_ net1382 vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09471__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17621_ clknet_leaf_111_wb_clk_i _03306_ _01562_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_95_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14833_ net1287 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17571__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11627__A1 _07588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17552_ clknet_leaf_13_wb_clk_i _03239_ _01535_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12101__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14764_ net1197 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__inv_2
XANTENNA__08087__A team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11976_ net2711 net234 net473 vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16503_ clknet_leaf_112_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[1\]
+ _00486_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13715_ net2782 _04102_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__nor2_1
XANTENNA__08518__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10927_ _06980_ _07227_ _07265_ _06921_ _07185_ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17483_ clknet_leaf_3_wb_clk_i _03170_ _01466_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14695_ net1346 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__inv_2
X_17963__1463 vssd1 vssd1 vccd1 vccd1 _17963__1463/HI net1463 sky130_fd_sc_hd__conb_1
XANTENNA__11940__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13646_ _03868_ _03880_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__xnor2_1
X_16434_ clknet_leaf_104_wb_clk_i _02188_ _00417_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10858_ _06158_ net374 net342 net341 net551 net539 vssd1 vssd1 vccd1 vccd1 _07198_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__14041__A2 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16365_ clknet_leaf_75_wb_clk_i net1634 _00348_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[88\]
+ sky130_fd_sc_hd__dfrtp_1
X_13577_ net984 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] _04022_ _04023_
+ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10789_ _04919_ _07125_ _07128_ vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18104_ net636 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_1
X_15316_ net1263 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12528_ net3048 net248 net405 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__mux2_1
X_16296_ clknet_leaf_73_wb_clk_i _02050_ _00279_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18035_ net1535 vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__buf_2
X_15247_ net1214 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12459_ net3024 net222 net413 vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__mux2_1
XANTENNA__13552__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16519__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15178_ net1272 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08550__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10366__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09220__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14129_ _04404_ _04411_ _04413_ _04414_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__or4_2
XFILLER_0_123_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout309 net313 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_2
XANTENNA__09084__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16669__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_77_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09670_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[22\] net959
+ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__and3_1
X_08621_ _04955_ _04957_ _04958_ _04960_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__or4_1
X_17819_ clknet_leaf_68_wb_clk_i net1630 _01759_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12011__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11618__A1 _07088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[19\] net893 vssd1
+ vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__and3_1
XANTENNA__10320__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08483_ net1087 net886 vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__and2_2
XANTENNA__11850__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10841__A2 _06636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14032__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09104_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[13\] net696 _05423_
+ _05424_ _05429_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11151__A _07449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09995__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16032__RESET_B _00026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09035_ _05338_ _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__nand2_1
XANTENNA__12681__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1231_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1329_A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16199__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13543__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold330 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[9\] vssd1 vssd1 vccd1 vccd1
+ net1946 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08460__A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold341 net124 vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold352 _02158_ vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout789_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold374 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[31\] vssd1 vssd1 vccd1 vccd1 net2001
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14099__A2 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold396 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 _04639_ vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__buf_4
Xfanout821 net824 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__buf_8
X_09937_ _06273_ _06274_ _06276_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__or3_1
XFILLER_0_102_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout832 team_01_WB.instance_to_wrap.cpu.RU0.next_ihit vssd1 vssd1 vccd1 vccd1 net832
+ sky130_fd_sc_hd__buf_1
Xfanout843 net846 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__buf_2
Xfanout854 net855 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_4
Xfanout865 net867 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__buf_2
XANTENNA__17594__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13806__A team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout876 team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1 vccd1
+ net876 sky130_fd_sc_hd__buf_2
XFILLER_0_99_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09868_ _06202_ _06203_ _06204_ _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__or4_1
Xfanout887 _04799_ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_8
Xhold1030 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[80\] vssd1 vssd1 vccd1 vccd1
+ net2646 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout898 net899 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1041 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ net1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[1\] net903 vssd1
+ vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__and3_1
Xhold1052 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[46\] vssd1 vssd1 vccd1 vccd1
+ net2668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2679 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[14\] net750 net744 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__a22o_1
Xhold1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1096 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2712 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11609__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11830_ net2699 net219 net487 vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__mux2_1
XANTENNA__10230__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09278__A2 _05615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11761_ net2264 net220 net497 vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__mux2_1
XANTENNA__11085__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12856__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11760__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13500_ net198 net194 _07826_ net644 vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10712_ _06934_ _07043_ _07051_ _06963_ _07048_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14480_ net1330 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__inv_2
XANTENNA__10832__A2 _06472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold701_A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11692_ _07808_ _07890_ vssd1 vssd1 vccd1 vccd1 _07891_ sky130_fd_sc_hd__nor2_1
XANTENNA__14023__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _03890_ _03891_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__or2_1
X_10643_ _06671_ _06707_ net543 vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10045__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09986__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16150_ clknet_leaf_96_wb_clk_i _01913_ _00138_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13362_ net585 _07684_ _03832_ _03831_ net564 vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__a32o_1
XANTENNA__11242__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10574_ _06910_ _06913_ vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__nor2_1
XANTENNA__10596__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09450__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15101_ net1262 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__inv_2
X_12313_ net1980 net251 net432 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16081_ clknet_leaf_103_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[3\]
+ _00069_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12591__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13293_ _03746_ _03778_ _04518_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15032_ net1171 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__inv_2
XANTENNA__13534__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12244_ net2635 net255 net439 vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__mux2_1
XANTENNA__08370__A team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_107_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_111_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08801__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12175_ net2944 net260 net449 vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__mux2_1
XANTENNA__16811__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11126_ net534 _06952_ _06954_ _07465_ net376 vssd1 vssd1 vccd1 vccd1 _07466_ sky130_fd_sc_hd__o311a_1
X_16983_ clknet_leaf_137_wb_clk_i _02670_ _00966_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11935__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15934_ net1394 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__inv_2
X_11057_ _07395_ _07396_ vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10008_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[1\] net823 net774 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__a22o_1
XANTENNA__09910__B1 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16961__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15865_ net1396 vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__inv_2
XANTENNA__09632__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17604_ clknet_leaf_71_wb_clk_i _03291_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14816_ net1243 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15796_ net1381 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__inv_2
XANTENNA__09269__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17535_ clknet_leaf_25_wb_clk_i _03222_ _01518_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14747_ net1308 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__inv_2
X_11959_ net575 _07945_ _07951_ vssd1 vssd1 vccd1 vccd1 _07952_ sky130_fd_sc_hd__and3_4
XFILLER_0_114_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17317__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11670__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10284__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17466_ clknet_leaf_45_wb_clk_i _03153_ _01449_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14678_ net1368 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16417_ clknet_leaf_79_wb_clk_i _02171_ _00400_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13629_ net982 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] _04066_ _04067_
+ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17397_ clknet_leaf_124_wb_clk_i _03084_ _01380_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09977__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16348_ clknet_leaf_78_wb_clk_i _02102_ _00331_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17467__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16279_ clknet_leaf_64_wb_clk_i _02033_ _00262_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13525__A1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18018_ net1518 vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_114_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11536__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08711__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16491__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10315__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12006__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07983_ team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 _04481_
+ sky130_fd_sc_hd__inv_2
XANTENNA__11845__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09722_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[21\] net807 net768 _06060_
+ _06061_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09901__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[23\] net753 _05991_
+ _05992_ net768 vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09542__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout272_A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\] net704 _04931_ _04943_
+ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_2_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09584_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[25\] net808 _05903_
+ _05906_ _05909_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08535_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[18\] net665 _04852_
+ _04858_ _04866_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12676__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10985__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1181_A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1279_A net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08466_ net1011 net891 vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__and2_2
XFILLER_0_37_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14005__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09680__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18033__1533 vssd1 vssd1 vccd1 vccd1 _18033__1533/HI net1533 sky130_fd_sc_hd__conb_1
XFILLER_0_50_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout704_A _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] net714 net710 vssd1 vssd1
+ vccd1 vccd1 _04737_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09968__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09432__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16834__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09018_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[9\] net895 vssd1
+ vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13516__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09286__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10290_ net1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[19\] net962
+ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11527__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12724__C1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 _01967_ vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _03532_ vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 net1798
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17962__1462 vssd1 vssd1 vccd1 vccd1 _17962__1462/HI net1462 sky130_fd_sc_hd__conb_1
Xhold193 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[1\] vssd1 vssd1 vccd1 vccd1
+ net1809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout640 net642 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11755__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout651 net652 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__buf_6
Xfanout662 _04811_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__buf_6
X_13980_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[48\] _04236_ _04259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__a22o_1
Xfanout673 net674 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__clkbuf_8
Xfanout684 _04783_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_8
Xfanout695 net696 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_8
X_12931_ _05453_ _07757_ _03694_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__o21ai_2
XANTENNA__13255__B team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16214__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12862_ net2503 net305 net381 vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
X_15650_ net1264 vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11813_ net2631 net254 net493 vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__mux2_1
X_14601_ net1377 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__inv_2
X_15581_ net1252 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__inv_2
XANTENNA__12586__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12793_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] net1056 net365 _03623_
+ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14532_ net1392 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__inv_2
X_17320_ clknet_leaf_22_wb_clk_i _03007_ _01303_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11744_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[3\] net718 net615 vssd1 vssd1
+ vccd1 vccd1 _07933_ sky130_fd_sc_hd__o21a_1
XANTENNA__10805__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16364__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17251_ clknet_leaf_21_wb_clk_i _02938_ _01234_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14463_ net1361 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13204__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11675_ net2680 net269 net499 vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09959__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13414_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] _05224_ vssd1 vssd1 vccd1
+ vccd1 _03875_ sky130_fd_sc_hd__xnor2_1
X_16202_ clknet_leaf_113_wb_clk_i _01962_ _00190_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17182_ clknet_leaf_48_wb_clk_i _02869_ _01165_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10626_ net553 _06965_ vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14394_ net1309 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__inv_2
XANTENNA__09423__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16133_ clknet_leaf_93_wb_clk_i _00024_ _00121_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_106_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13345_ _04482_ _07678_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__nand2_1
X_10557_ net545 net536 _06858_ vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__or3_1
XFILLER_0_52_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09974__A3 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13507__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16064_ clknet_leaf_121_wb_clk_i _01857_ _00052_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09196__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13276_ net1656 net825 _07650_ _03765_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10488_ _06750_ _06819_ _06823_ _06827_ _05902_ vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_27_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15015_ net1301 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12227_ net2780 net224 net439 vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__mux2_1
XANTENNA__15926__A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12158_ net3026 net190 net447 vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__mux2_1
XANTENNA__11665__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ net345 _06409_ _07439_ _07448_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__o31a_2
XFILLER_0_97_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16966_ clknet_leaf_40_wb_clk_i _02653_ _00949_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12089_ net3184 net317 net462 vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__mux2_1
X_15917_ net1411 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11297__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16897_ clknet_leaf_48_wb_clk_i _02584_ _00880_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15661__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15848_ net1363 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12496__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15779_ net1307 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08320_ net1146 net1154 net1151 net1149 vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_115_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12797__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17518_ clknet_leaf_5_wb_clk_i _03205_ _01501_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08706__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08251_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[30\] net1779 net1037 vssd1 vssd1
+ vccd1 vccd1 _03436_ sky130_fd_sc_hd__mux2_1
X_17449_ clknet_leaf_10_wb_clk_i _03136_ _01432_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16857__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08182_ net2586 net2351 net1053 vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08622__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10980__A1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09537__C net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08441__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10980__B2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1027_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16237__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_A _07947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09705_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[21\] net945 vssd1
+ vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout654_A _04819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1396_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09636_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[23\] net975
+ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__and3_1
XANTENNA__16387__CLK clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17632__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09567_ _04491_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[25\] net965 vssd1
+ vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout821_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout919_A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11604__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[18\] net882 vssd1
+ vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09498_ _04706_ _05836_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09653__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08449_ net1083 net896 vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__and2_2
XFILLER_0_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11323__B team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ net1155 _04713_ net720 _04751_ vssd1 vssd1 vccd1 vccd1 _07756_ sky130_fd_sc_hd__o22a_2
XFILLER_0_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09405__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10411_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[27\] net954
+ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08613__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11391_ team_01_WB.instance_to_wrap.cpu.f0.i\[30\] _07716_ _07717_ vssd1 vssd1 vccd1
+ vccd1 _03393_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13030__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13130_ net2391 net847 net632 team_01_WB.instance_to_wrap.a1.ADR_I\[13\] vssd1 vssd1
+ vccd1 vccd1 _02011_ sky130_fd_sc_hd__a22o_1
XANTENNA__17012__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10342_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[17\] net962
+ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10971__A1 _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10971__B2 _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13061_ net3172 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[33\] net866 vssd1 vssd1
+ vccd1 vccd1 _02064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10273_ net1120 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[19\] net953
+ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12012_ net2161 net289 net470 vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1402 net1404 vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__buf_4
XANTENNA_input48_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1413 net1414 vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__buf_2
XFILLER_0_40_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_126_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13266__A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17162__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16820_ clknet_leaf_12_wb_clk_i _02507_ _00803_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_54_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout470 _07953_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_50_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout481 _07949_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16751_ clknet_leaf_142_wb_clk_i _02438_ _00734_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout492 _07944_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13963_ _04231_ _04237_ _04239_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_31_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13673__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09341__A1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15702_ net1201 vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__inv_2
X_12914_ net362 _03684_ net1025 vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__o21ai_2
X_13894_ _04140_ net571 _04198_ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__and3_1
X_16682_ clknet_leaf_2_wb_clk_i _02369_ _00665_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15633_ net1288 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__inv_2
X_12845_ net3053 net271 net380 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__mux2_1
XANTENNA__13425__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10239__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ net1028 _07231_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15564_ net1197 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09644__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17303_ clknet_leaf_138_wb_clk_i _02990_ _01286_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08526__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14515_ net1407 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11727_ net721 _07323_ net615 _07918_ vssd1 vssd1 vccd1 vccd1 _07919_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15495_ net1327 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17234_ clknet_leaf_134_wb_clk_i _02921_ _01217_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11658_ net721 _07171_ net616 _07863_ vssd1 vssd1 vccd1 vccd1 _07864_ sky130_fd_sc_hd__o211a_1
X_14446_ net1400 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11739__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10609_ _06438_ net373 net546 vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__mux2_1
X_14377_ net1318 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__inv_2
X_17165_ clknet_leaf_138_wb_clk_i _02852_ _01148_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11589_ _07805_ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold907 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold918 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[112\] vssd1 vssd1 vccd1 vccd1
+ net2534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16116_ clknet_leaf_101_wb_clk_i _01891_ _00104_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13328_ team_01_WB.instance_to_wrap.cpu.f0.i\[16\] _03743_ _03801_ net586 vssd1 vssd1
+ vccd1 vccd1 _03806_ sky130_fd_sc_hd__o211a_1
XANTENNA__12951__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17096_ clknet_leaf_24_wb_clk_i _02783_ _01079_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold929 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16047_ clknet_leaf_87_wb_clk_i _01840_ _00035_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_13259_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] net1063 _07710_ vssd1 vssd1 vccd1
+ vccd1 _03751_ sky130_fd_sc_hd__or3_1
XANTENNA__17505__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18032__1532 vssd1 vssd1 vccd1 vccd1 _18032__1532/HI net1532 sky130_fd_sc_hd__conb_1
Xhold1607 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17998_ net1498 vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_hd__buf_2
Xhold1618 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net3234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1629 team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 net3245
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09092__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16949_ clknet_leaf_121_wb_clk_i _02636_ _00932_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13664__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10031__C net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09421_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[28\] net657 net653 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09352_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[25\] net661 net657 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[25\]
+ _05684_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__a221o_1
XANTENNA__08209__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08303_ net989 net967 vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_118_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17961__1461 vssd1 vssd1 vccd1 vccd1 _17961__1461/HI net1461 sky130_fd_sc_hd__conb_1
XFILLER_0_74_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09283_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[22\] net919
+ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_60_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12954__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10650__A0 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08234_ net2003 net2837 net1047 vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13195__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08165_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[116\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[108\]
+ net1040 vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout402_A _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1144_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08096_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[28\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[31\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[30\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17185__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1311_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1409_A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10206__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09564__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout771_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ _05303_ _05337_ net603 vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_3_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17906__1426 vssd1 vssd1 vccd1 vccd1 _17906__1426/HI net1426 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_86_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10960_ _07117_ _07199_ net514 vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11130__A1 _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11130__B2 _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09874__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09619_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[24\] net737 _05939_ _05946_
+ _05947_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09730__C net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11681__A2 _07611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ net562 _07208_ _07209_ _07230_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__a31oi_4
X_12630_ net2960 net208 net391 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14080__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[26\] net250 net401 vssd1
+ vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12864__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11433__A2 _07701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14300_ net1355 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__inv_2
X_11512_ net1648 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\] net877 vssd1 vssd1
+ vccd1 vccd1 _03337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15280_ net1224 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__inv_2
X_12492_ net2540 net222 net409 vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14231_ net1636 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13186__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11443_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] team_01_WB.instance_to_wrap.cpu.f0.i\[3\]
+ _07673_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1 _07746_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14162_ _04188_ _04441_ _04195_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__o21a_1
XANTENNA__12933__A2 _03697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11374_ _04478_ _07702_ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09177__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10944__A1 _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13113_ net1732 net843 net635 team_01_WB.instance_to_wrap.a1.ADR_I\[30\] vssd1 vssd1
+ vccd1 vccd1 _02028_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10325_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[18\] net945 vssd1
+ vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_128_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14093_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] _04249_ _04265_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\]
+ _04379_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ net1609 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
X_13044_ net2409 net2300 net857 vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__mux2_1
XANTENNA__09474__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10256_ _06594_ _06595_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__nand2b_1
XANTENNA__16552__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1210 net1211 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1221 net1227 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1232 net1235 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__buf_4
X_17852_ clknet_leaf_65_wb_clk_i net2350 _01792_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12104__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ _06526_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__inv_2
XANTENNA__10413__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10172__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1243 net1245 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1254 net1257 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__buf_4
XFILLER_0_94_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16803_ clknet_leaf_21_wb_clk_i _02490_ _00786_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1265 net1269 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__clkbuf_2
Xfanout1276 net1277 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__buf_4
X_17783_ clknet_leaf_62_wb_clk_i _03459_ _01723_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[53\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout1287 net1294 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__buf_4
X_14995_ net1280 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1298 net1302 vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11943__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09314__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16734_ clknet_leaf_48_wb_clk_i _02421_ _00717_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13946_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__or2_4
XANTENNA__09865__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16665_ clknet_leaf_47_wb_clk_i _02352_ _00648_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09640__C net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11672__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13877_ team_01_WB.EN_VAL_REG net2667 vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__and2b_1
X_15616_ net1243 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__inv_2
XANTENNA__10880__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12828_ net3247 net640 net607 _03648_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14071__B1 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16596_ clknet_leaf_127_wb_clk_i _02283_ _00579_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_130_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15547_ net1183 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12759_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] net1054 net363 _03600_
+ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15478_ net1224 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17217_ clknet_leaf_42_wb_clk_i _02904_ _01200_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14429_ net1365 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12924__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17148_ clknet_leaf_37_wb_clk_i _02835_ _01131_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold704 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09087__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold715 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold737 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[25\] vssd1 vssd1 vccd1 vccd1
+ net2353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09970_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[3\] net780 net771 _06293_
+ _06298_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__a2111o_1
Xhold748 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
X_17079_ clknet_leaf_138_wb_clk_i _02766_ _01062_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08921_ net603 _05258_ _05259_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_21_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08356__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[3\] net903 vssd1
+ vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__and3_1
XANTENNA__12014__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1404 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3020 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10163__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1415 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1426 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08783_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[0\] net881 vssd1
+ vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__and3_1
Xhold1437 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1448 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[59\] vssd1 vssd1 vccd1 vccd1
+ net3064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout185_A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1459 team_01_WB.instance_to_wrap.cpu.f0.num\[18\] vssd1 vssd1 vccd1 vccd1 net3075
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11853__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09856__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12860__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1094_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11154__A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08447__B net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09404_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[27\] net670 net650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[27\]
+ _05743_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__a221o_1
XANTENNA__10871__A0 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14062__B1 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[24\] net661 net651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[24\]
+ _05664_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12684__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16425__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_830 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1261_A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10623__B1 _06921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1359_A net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09266_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[20\] net672 net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__a22o_1
XANTENNA__09559__A _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13168__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08217_ net2969 net2717 net1049 vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__mux2_1
XANTENNA__11601__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09197_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[17\] net931 vssd1
+ vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_75_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08148_ _04583_ _04599_ _04616_ _04617_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__and4bb_1
XANTENNA__09241__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08044__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout986_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08079_ net1814 net569 _04525_ _04553_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__a22o_1
X_10110_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[6\] net774 net771 vssd1
+ vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11090_ _04706_ _05835_ _06883_ _07428_ _07429_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__o311a_1
XFILLER_0_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[0\] net948 vssd1
+ vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__and3_1
Xhold20 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10154__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[2\] vssd1 vssd1 vccd1 vccd1
+ net1647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold42 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[24\] vssd1 vssd1 vccd1 vccd1
+ net1658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 team_01_WB.instance_to_wrap.cpu.f0.write_data\[28\] vssd1 vssd1 vccd1 vccd1
+ net1669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[105\] vssd1 vssd1 vccd1 vccd1
+ net1680 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12859__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13628__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold75 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[4\] vssd1 vssd1 vccd1 vccd1 net1691
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11763__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13800_ _01835_ _04176_ _04180_ _04159_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__o22a_1
Xhold86 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[10\] vssd1 vssd1 vccd1 vccd1
+ net1702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 _02014_ vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ net1176 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__inv_2
X_11992_ net575 _07793_ _07951_ vssd1 vssd1 vccd1 vccd1 _07953_ sky130_fd_sc_hd__and3_1
XANTENNA__09847__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10943_ _07156_ _07282_ net515 vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__mux2_1
X_13731_ team_01_WB.instance_to_wrap.a1.WRITE_I _04508_ team_01_WB.instance_to_wrap.a1.curr_state\[0\]
+ _04509_ net3153 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10862__A0 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16450_ clknet_leaf_21_wb_clk_i _02204_ _00433_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13662_ net199 net195 _04501_ net645 vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10874_ _05898_ net504 _06811_ _05931_ net548 net538 vssd1 vssd1 vccd1 vccd1 _07214_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15401_ net1229 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12613_ net3261 net279 net396 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16381_ clknet_leaf_76_wb_clk_i net2737 _00364_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12594__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13593_ _03903_ _04030_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12603__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12544_ net2932 net251 net404 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__mux2_1
X_15332_ net1238 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09480__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08373__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18031__1531 vssd1 vssd1 vccd1 vccd1 _18031__1531/HI net1531 sky130_fd_sc_hd__conb_1
XFILLER_0_87_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16918__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18051_ net1551 vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__buf_2
XFILLER_0_35_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12475_ net2197 net257 net411 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__mux2_1
X_15263_ net1254 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17002_ clknet_leaf_2_wb_clk_i _02689_ _00985_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12906__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13564__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14214_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] vssd1 vssd1 vccd1
+ vccd1 _02273_ sky130_fd_sc_hd__clkbuf_1
X_11426_ _07681_ _07700_ vssd1 vssd1 vccd1 vccd1 _07738_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_6 _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08035__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09232__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15194_ net1190 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_54_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_39_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14145_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[15\] _04253_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[63\]
+ _04429_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__a221o_1
XANTENNA__11938__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ net1065 _07677_ vssd1 vssd1 vccd1 vccd1 _07686_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10393__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10308_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[18\] net971
+ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__and3_1
X_14076_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[92\] _04241_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[28\]
+ _04363_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__a221o_1
X_11288_ _04734_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] net1155 vssd1 vssd1
+ vccd1 vccd1 _07628_ sky130_fd_sc_hd__or3b_1
XANTENNA__09635__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13027_ net2091 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[67\] net864 vssd1 vssd1
+ vccd1 vccd1 _02098_ sky130_fd_sc_hd__mux2_1
X_17904_ net1424 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_0_24_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10239_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[9\] net820 net806 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_89_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17960__1460 vssd1 vssd1 vccd1 vccd1 _17960__1460/HI net1460 sky130_fd_sc_hd__conb_1
Xfanout1040 net1045 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__buf_2
Xfanout1051 net1053 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__clkbuf_4
X_17835_ clknet_leaf_71_wb_clk_i _03511_ _01775_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[105\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1062 team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 net1062
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1073 net1075 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1084 net1086 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__buf_2
Xfanout1095 net1096 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__buf_2
XANTENNA__13454__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17766_ clknet_leaf_56_wb_clk_i _03442_ _01706_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_83_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08548__A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14978_ net1312 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16717_ clknet_leaf_139_wb_clk_i _02404_ _00700_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13929_ _04217_ _04219_ _04220_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__and3_4
XFILLER_0_92_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16448__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17697_ clknet_leaf_101_wb_clk_i _03381_ _01638_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16648_ clknet_leaf_22_wb_clk_i _02335_ _00631_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14044__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16579_ clknet_leaf_19_wb_clk_i _02266_ _00562_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09120_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[14\] net921 vssd1
+ vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11702__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16598__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17843__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08714__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09051_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[12\] net937 vssd1
+ vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17905__1425 vssd1 vssd1 vccd1 vccd1 _17905__1425/HI net1425 sky130_fd_sc_hd__conb_1
XFILLER_0_60_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12009__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08002_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1 vccd1 vccd1
+ _04500_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold501 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11848__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold523 team_01_WB.instance_to_wrap.cpu.f0.num\[24\] vssd1 vssd1 vccd1 vccd1 net2139
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13570__A2 _07251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold545 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold556 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10384__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold567 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09953_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[3\] net813 net759 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__a22o_1
Xhold589 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
X_08904_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[2\] net921 vssd1
+ vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__and3_1
XANTENNA__15844__A net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ net1134 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[5\] net954 vssd1
+ vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__and3_1
XANTENNA__10136__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1107_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1201 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[90\] vssd1 vssd1 vccd1 vccd1
+ net2817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 _03509_ vssd1 vssd1 vccd1 vccd1 net2828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17223__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08835_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[1\] net690 net660 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__a22o_1
Xhold1223 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2839 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1234 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 net2850
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12679__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1245 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2861 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout567_A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1256 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2872 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13364__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[4\] net700 _05088_ _05092_
+ _05094_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__a2111o_1
Xhold1267 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2894 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09829__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1289 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08697_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[7\] net700 _05007_ _05025_
+ net706 vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__a2111o_1
XANTENNA__17373__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13811__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout901_A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09318_ _05657_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10590_ _06897_ _06929_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__or2_1
XANTENNA__09462__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09249_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[21\] net689 net660 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[21\]
+ _05588_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13546__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12260_ net2908 net224 net435 vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11211_ net530 _07503_ _07549_ _07070_ vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_101_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08568__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10662__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ net2127 net191 net445 vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__mux2_1
XANTENNA__13561__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11142_ _05262_ net339 _07014_ _07481_ vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__a31o_1
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
XFILLER_0_25_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XANTENNA__13313__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15950_ net1391 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__inv_2
X_11073_ _05566_ _06707_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__or2_1
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
X_10024_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[1\] net777 _06362_ _06363_
+ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14901_ net1221 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15881_ net1383 vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__inv_2
XANTENNA__12589__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17620_ clknet_leaf_110_wb_clk_i _03305_ _01561_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13274__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14832_ net1270 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__inv_2
XANTENNA__17716__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17551_ clknet_leaf_141_wb_clk_i _03238_ _01534_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_101_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14763_ net1327 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12824__A1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11975_ net2237 net265 net472 vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__mux2_1
XANTENNA__12824__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16502_ clknet_leaf_108_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[0\]
+ _00485_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13714_ _04102_ _04119_ _04126_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[5\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_135_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10926_ _06980_ _07227_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__nor2_1
X_17482_ clknet_leaf_2_wb_clk_i _03169_ _01465_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14026__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14694_ net1343 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16740__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16433_ clknet_leaf_104_wb_clk_i _02187_ _00416_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10857_ net371 _07195_ _07196_ net341 _04970_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__o32a_1
XFILLER_0_39_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13645_ net983 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] _04079_ _04080_
+ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08815__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16364_ clknet_leaf_78_wb_clk_i _02118_ _00347_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_140_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09453__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13576_ net729 _07231_ net984 vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__a21oi_1
X_10788_ net336 _07127_ _07126_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18103_ net638 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15315_ net1234 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12527_ net3165 net215 net405 vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__mux2_1
X_16295_ clknet_leaf_65_wb_clk_i _02049_ _00278_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16890__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18034_ net1534 vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__buf_2
XFILLER_0_125_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15246_ net1285 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__inv_2
XANTENNA__08831__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12458_ net2963 net225 net411 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08559__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11409_ _07701_ _07711_ _07727_ net325 vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__o211a_1
XANTENNA__13552__A2 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15177_ net1229 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__inv_2
X_12389_ net2611 net293 net425 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10366__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12760__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16120__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17246__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14128_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[86\] _04245_ _04396_ _04152_
+ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14059_ _04347_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__inv_2
XANTENNA__10118__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12499__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08620_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[11\] net667 net655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[11\]
+ _04959_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__a221o_1
XANTENNA__17396__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08731__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17818_ clknet_leaf_85_wb_clk_i _03494_ _01758_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08709__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08551_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[19\] net889
+ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__and3_1
X_17749_ clknet_leaf_73_wb_clk_i _03425_ _01689_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10826__A0 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08482_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[23\] net882 vssd1
+ vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09692__B1 _06030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10841__A3 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08217__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09103_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[13\] net690 _05431_
+ _05433_ _05440_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_94_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11151__B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08444__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12962__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout315_A _07939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09034_ _05339_ _05373_ net602 vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__mux2_4
XANTENNA__13528__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1057_A team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08741__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold320 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1
+ net1936 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13543__A2 _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold331 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08460__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1224_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[4\] vssd1 vssd1 vccd1 vccd1
+ net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold375 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout800 _04646_ vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_8
Xhold386 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold397 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 net814 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__buf_6
XFILLER_0_99_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09936_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[4\] net811 net798 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[4\]
+ _06275_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__a221o_1
Xfanout822 net824 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__buf_6
XANTENNA__16613__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10109__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11306__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout833 net834 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout844 net846 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__buf_2
Xfanout855 net856 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__buf_2
Xfanout866 net867 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09572__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout851_A _03731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[12\] net741 _06205_ _06206_
+ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__a211o_1
Xfanout877 team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1 vccd1
+ net877 sky130_fd_sc_hd__clkbuf_4
Xfanout888 net891 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__buf_4
Xhold1020 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[15\] vssd1 vssd1 vccd1 vccd1 net2636
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout899 _04788_ vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__buf_4
XANTENNA_fanout949_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18030__1530 vssd1 vssd1 vccd1 vccd1 _18030__1530/HI net1530 sky130_fd_sc_hd__conb_1
Xhold1042 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[27\] vssd1 vssd1 vccd1 vccd1
+ net2658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08818_ net1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[1\] net880 vssd1
+ vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1053 _03452_ vssd1 vssd1 vccd1 vccd1 net2669 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12202__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09798_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[14\] net789 net741 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__a22o_1
Xhold1064 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1075 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[48\] vssd1 vssd1 vccd1 vccd1
+ net2691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2702 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16763__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2713 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[4\] net925 vssd1
+ vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12806__B2 _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14918__A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10817__A0 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11760_ net2995 net223 net495 vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__mux2_1
XANTENNA__14008__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09683__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ net554 _07050_ vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11691_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _07805_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\]
+ vssd1 vssd1 vccd1 vccd1 _07890_ sky130_fd_sc_hd__a21oi_1
XANTENNA__17119__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11342__A team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10642_ net375 net372 net549 vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__mux2_1
X_13430_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] net595 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\]
+ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09435__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ _04484_ _07683_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10573_ _04741_ _04743_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__or2_1
X_15100_ net1174 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12312_ net2772 net227 net432 vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16080_ clknet_leaf_103_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[2\]
+ _00068_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[2\] sky130_fd_sc_hd__dfrtp_1
X_13292_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] _03744_ vssd1 vssd1 vccd1 vccd1
+ _03778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12243_ net3000 net261 net441 vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15031_ net1200 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08370__B team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10979__S0 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12174_ net2988 net231 net448 vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__mux2_1
XANTENNA__09185__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11125_ net534 _07453_ vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__nand2_1
XANTENNA__08961__A2 _05300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16982_ clknet_leaf_1_wb_clk_i _02669_ _00965_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15933_ net1411 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__inv_2
X_11056_ net557 _06280_ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10007_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[1\] net820 net814 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__a22o_1
XANTENNA__09910__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12112__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15864_ net1385 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__inv_2
X_17904__1424 vssd1 vssd1 vccd1 vccd1 _17904__1424/HI net1424 sky130_fd_sc_hd__conb_1
XANTENNA__10520__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17603_ clknet_leaf_71_wb_clk_i _03290_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_14815_ net1254 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__inv_2
XANTENNA__08529__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15795_ net1381 vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__inv_2
XANTENNA__11951__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17534_ clknet_leaf_45_wb_clk_i _03221_ _01517_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14746_ net1310 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__inv_2
X_11958_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\]
+ vssd1 vssd1 vccd1 vccd1 _07951_ sky130_fd_sc_hd__and2b_2
XFILLER_0_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17465_ clknet_leaf_47_wb_clk_i _03152_ _01448_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10909_ _07100_ _07242_ _07248_ net329 _07247_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14677_ net1378 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__inv_2
X_11889_ net3188 net319 net486 vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16416_ clknet_leaf_106_wb_clk_i _02170_ _00399_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13628_ net723 _07269_ net1068 vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09426__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17396_ clknet_leaf_13_wb_clk_i _03083_ _01379_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13222__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16347_ clknet_leaf_86_wb_clk_i _02101_ _00330_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13559_ net185 _04007_ _04008_ net725 vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__a211o_1
XFILLER_0_125_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10587__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09657__A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16278_ clknet_leaf_67_wb_clk_i _02032_ _00261_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08561__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18017_ net1517 vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_57_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13525__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15229_ net1262 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11536__B2 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09095__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08952__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07982_ team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 _04480_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10034__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire917_A net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16786__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09721_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[21\] net756 _06043_ _06044_
+ _06046_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_59_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12022__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[23\] net782 _05970_ _05971_
+ _05977_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10511__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08603_ _04935_ _04936_ _04939_ _04942_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__or4_2
X_09583_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[25\] net822 net752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11861__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08534_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[18\] net649 _04848_
+ _04851_ _04857_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13997__C1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10985__B _06398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08465_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[23\] net882
+ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout432_A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1174_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13213__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09417__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08396_ _04733_ _04735_ _04734_ _04731_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_18_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17411__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12692__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1341_A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09567__A _04491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08471__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09017_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[9\] net880 vssd1
+ vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__and3_1
XANTENNA__08902__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13516__A2 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17561__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11527__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold150 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold161 net158 vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__C1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold183 net92 vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout630 _03738_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_4
Xfanout641 net642 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__buf_2
Xfanout652 _04821_ vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__buf_8
X_09919_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[4\] net785 net760 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__a22o_1
Xfanout663 _04808_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__buf_8
Xfanout674 _04794_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__buf_4
Xfanout685 _04780_ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_8
Xfanout696 _04768_ vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__buf_8
X_12930_ net359 _03695_ _03696_ net872 net3191 vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_124_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10502__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08349__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12861_ net2181 net309 net382 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11771__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14600_ net1339 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__inv_2
X_11812_ net2760 net230 net494 vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15580_ net1174 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
XANTENNA__09656__B1 _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12792_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[12\] _07520_ net1028 vssd1 vssd1
+ vccd1 vccd1 _03623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14531_ net1408 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__inv_2
X_11743_ net719 net322 vssd1 vssd1 vccd1 vccd1 _07932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17250_ clknet_leaf_32_wb_clk_i _02937_ _01233_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09408__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13204__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14462_ net1360 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17091__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11674_ _07874_ _07876_ net614 vssd1 vssd1 vccd1 vccd1 _07877_ sky130_fd_sc_hd__mux2_2
X_16201_ clknet_leaf_113_wb_clk_i _01961_ _00189_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13413_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _05116_ _07641_ _07640_
+ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17181_ clknet_leaf_21_wb_clk_i _02868_ _01164_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10625_ net529 net503 vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14393_ net1309 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__inv_2
XANTENNA__16659__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12963__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16132_ clknet_leaf_93_wb_clk_i _00023_ _00120_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13344_ net1894 net827 _03816_ _03818_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__o22a_1
X_10556_ net545 _05899_ _06895_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__a21o_1
XFILLER_0_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10974__C1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16063_ clknet_leaf_121_wb_clk_i _01856_ _00051_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10416__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13275_ net586 _03763_ _03764_ net565 vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__a22o_1
X_10487_ _05869_ _05870_ vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__or2_1
XANTENNA__12107__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11518__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15014_ net1295 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__inv_2
X_12226_ net3179 net191 net439 vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11946__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12157_ _07791_ net576 _07942_ vssd1 vssd1 vccd1 vccd1 _07958_ sky130_fd_sc_hd__and3_4
XFILLER_0_20_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11108_ _07071_ _07447_ _07444_ _07441_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__o211a_1
X_12088_ net3260 net319 net462 vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__mux2_1
X_16965_ clknet_leaf_40_wb_clk_i _02652_ _00948_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16039__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13140__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11039_ _07259_ _07373_ _07377_ _07378_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__and4b_1
X_15916_ net1398 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__inv_2
XANTENNA__09895__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16896_ clknet_leaf_30_wb_clk_i _02583_ _00879_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15847_ net1351 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16189__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09647__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15778_ net1306 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08556__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09151__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09111__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17517_ clknet_leaf_140_wb_clk_i _03204_ _01500_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13181__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14729_ net1344 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08250_ net3088 net3015 net1047 vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__mux2_1
X_17448_ clknet_leaf_22_wb_clk_i _03135_ _01431_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08181_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[100\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[92\]
+ net1039 vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ clknet_leaf_22_wb_clk_i _03066_ _01362_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12954__A0 team_01_WB.instance_to_wrap.cpu.f0.write_data\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_9_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_65_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08722__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12017__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10326__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09178__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11856__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_74_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13131__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ net1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[21\] net953
+ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09635_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[23\] net943
+ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__and3_1
XANTENNA__09350__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14468__A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1291_A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A _04825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1389_A net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09566_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[25\] net968
+ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__and3_1
XANTENNA__08466__A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11604__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[18\] net919
+ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__and3_1
XANTENNA__11445__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13985__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09497_ _04706_ _05836_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08448_ net1109 net1112 net1114 net1106 vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__and4b_1
XFILLER_0_33_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_83_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13198__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08379_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\]
+ net1156 vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__and3b_1
XFILLER_0_68_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11748__A1 _07489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12945__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10410_ _06748_ _06749_ _05934_ _05967_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_22_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11390_ _07717_ _07718_ _04465_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__mux2_1
XANTENNA__09810__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08632__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17903__1423 vssd1 vssd1 vccd1 vccd1 _17903__1423/HI net1423 sky130_fd_sc_hd__conb_1
X_10341_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[17\] net953 vssd1
+ vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__and3_1
X_13060_ net2715 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[34\] net858 vssd1 vssd1
+ vccd1 vccd1 _02065_ sky130_fd_sc_hd__mux2_1
XANTENNA__09169__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10272_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[19\] net740 _06609_ _06610_
+ _06611_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__a2111o_1
X_12011_ net2693 net257 net468 vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__mux2_1
XANTENNA__11766__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08916__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13370__B1 _07650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17307__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1403 net1404 vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__buf_4
Xfanout1414 net1415 vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_92_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout460 _07955_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13122__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout471 _07952_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_50_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout482 _07949_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_4
XFILLER_0_45_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16750_ clknet_leaf_3_wb_clk_i _02437_ _00733_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13962_ _04218_ _04242_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__nor2_4
Xfanout493 _07944_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11133__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13673__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17457__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15701_ net1223 vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_79_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12913_ _04881_ net578 vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__nor2_1
XANTENNA__09341__A2 _05678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12597__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16681_ clknet_leaf_8_wb_clk_i _02368_ _00664_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13893_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _04198_
+ sky130_fd_sc_hd__a21o_1
X_15632_ net1224 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__inv_2
X_12844_ net2010 net245 net379 vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08807__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15563_ net1295 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12775_ net1865 net641 net608 _03611_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16481__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17302_ clknet_leaf_2_wb_clk_i _02989_ _01285_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14514_ net1394 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[6\] net718 vssd1 vssd1 vccd1
+ vccd1 _07918_ sky130_fd_sc_hd__or2_1
X_15494_ net1324 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13189__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17233_ clknet_leaf_14_wb_clk_i _02920_ _01216_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14445_ net1378 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__inv_2
X_11657_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[20\] net715 vssd1 vssd1 vccd1
+ vccd1 _07863_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11739__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12936__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10608_ _06946_ _06947_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__nor2_1
X_17164_ clknet_leaf_134_wb_clk_i _02851_ _01147_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14376_ net1318 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09638__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11588_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] _07803_ vssd1 vssd1
+ vccd1 vccd1 _07805_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16115_ clknet_leaf_101_wb_clk_i _01890_ _00103_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold908 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
X_13327_ net1678 net826 _03805_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__o21a_1
Xhold919 _02143_ vssd1 vssd1 vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[31\] net689 net670 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17095_ clknet_leaf_16_wb_clk_i _02782_ _01078_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16046_ clknet_leaf_107_wb_clk_i _01839_ _00034_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
X_13258_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] _03749_ vssd1 vssd1 vccd1 vccd1
+ _03750_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11676__S net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ net2686 net257 net443 vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10175__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13189_ net20 net837 net630 net2233 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09580__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17997_ net1497 vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__buf_2
Xhold1608 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1619 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3235 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_109_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13113__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15672__A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16948_ clknet_leaf_13_wb_clk_i _02635_ _00931_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13664__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09670__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16879_ clknet_leaf_142_wb_clk_i _02566_ _00862_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_09420_ net560 _05759_ _05737_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12300__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08717__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11427__B1 _07699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11424__B _07701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09351_ _05689_ _05690_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08302_ net1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[30\] net966
+ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_118_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09282_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[22\] net934
+ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_118_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ net2691 net2560 net1046 vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10650__A1 _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout228_A _07900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11440__A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08164_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[117\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[109\]
+ net1039 vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__mux2_1
XANTENNA__09399__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08225__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08452__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16204__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08095_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[25\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[24\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[27\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__or4_1
XANTENNA__15847__A net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1137_A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14144__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10166__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11902__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16354__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] net703 _05320_ _05336_
+ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA_fanout764_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09859__B1 _04678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09323__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout931_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11615__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09618_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[24\] net796 net776 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__a22o_1
XANTENNA__12210__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10890_ _07054_ _07228_ _07229_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09549_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[28\] net801 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[28\]
+ _05884_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11053__C net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12560_ net3218 net213 net401 vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08924__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11511_ net1816 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] net877 vssd1 vssd1
+ vccd1 vccd1 _03338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12491_ net1925 net225 net407 vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__mux2_1
XANTENNA__12918__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14230_ net2400 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_24_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_126_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11442_ _07676_ _07745_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__nor2_1
XANTENNA__08598__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11197__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13591__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14161_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[3\] _04187_ vssd1 vssd1 vccd1
+ vccd1 _04441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11373_ team_01_WB.instance_to_wrap.cpu.f0.i\[15\] _07682_ vssd1 vssd1 vccd1 vccd1
+ _07702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10944__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13112_ net1742 net844 net631 team_01_WB.instance_to_wrap.a1.ADR_I\[31\] vssd1 vssd1
+ vccd1 vccd1 _02029_ sky130_fd_sc_hd__a22o_1
X_10324_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[18\] net957
+ vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__and3_1
XANTENNA_input60_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14135__A2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14092_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[29\] _04267_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[77\]
+ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13277__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13343__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17920_ net1608 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
X_13043_ net2574 net2368 net864 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__mux2_1
X_10255_ net340 _06593_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1200 net1202 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__clkbuf_4
Xfanout1211 net1236 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__buf_2
X_17851_ clknet_leaf_68_wb_clk_i net1877 _01791_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10186_ net627 _06525_ _06502_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__o21ai_4
Xfanout1222 net1227 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_33_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09193__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1233 net1235 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1244 net1245 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__clkbuf_4
X_16802_ clknet_leaf_35_wb_clk_i _02489_ _00785_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1255 net1257 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16847__CLK clknet_leaf_143_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17782_ clknet_leaf_56_wb_clk_i _03458_ _01722_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[52\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout1266 net1268 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__buf_4
X_14994_ net1233 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__inv_2
Xfanout1277 net1303 vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__buf_2
Xfanout1288 net1294 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__buf_4
Xfanout290 _07896_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_2
Xfanout1299 net1301 vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__buf_4
X_16733_ clknet_leaf_20_wb_clk_i _02420_ _00716_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09314__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13945_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__nor2_2
XFILLER_0_117_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16664_ clknet_leaf_28_wb_clk_i _02351_ _00647_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12120__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13876_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\] _04186_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.lcd_en sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11672__A3 _07809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16997__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15615_ net1244 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__inv_2
X_12827_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] net1057 net366 _03647_
+ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__a22o_1
XANTENNA__09078__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16595_ clknet_leaf_117_wb_clk_i _02282_ _00578_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_56_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15546_ net1192 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12758_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[23\] _07111_ net1026 vssd1 vssd1
+ vccd1 vccd1 _03600_ sky130_fd_sc_hd__mux2_1
XANTENNA__08834__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10632__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11709_ net2342 net253 net501 vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16227__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15477_ net1223 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12689_ net1924 net225 net383 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17216_ clknet_leaf_29_wb_clk_i _02903_ _01199_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14428_ net1365 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08589__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_96_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15667__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17147_ clknet_leaf_17_wb_clk_i _02834_ _01130_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13582__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold705 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14359_ net1350 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__inv_2
Xhold716 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold727 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 net2343
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10307__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14126__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16377__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09665__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17078_ clknet_leaf_141_wb_clk_i _02765_ _01061_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17622__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08920_ net603 _05258_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__a21o_1
X_16029_ net1351 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10148__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08851_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[3\] net908 vssd1
+ vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1405 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1427 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net3043 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17772__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08782_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[0\] net892 vssd1
+ vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__and3_1
Xhold1438 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3054 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13637__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10042__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1449 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3065 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09305__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11112__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12030__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17902__1422 vssd1 vssd1 vccd1 vccd1 _17902__1422/HI net1422 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_81_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17002__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09403_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[27\] net904
+ net664 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[27\] vssd1 vssd1 vccd1
+ vccd1 _05743_ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10871__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout345_A _04748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1087_A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[24\] net695 _05673_
+ net707 vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08744__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09265_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[20\] net687 net686 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[20\]
+ _05597_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout512_A _05931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1254_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08216_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[65\] net2068 net1050 vssd1 vssd1
+ vccd1 vccd1 _03471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09196_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[17\] net893 vssd1
+ vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11179__A2 _07065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08147_ _04465_ team_01_WB.instance_to_wrap.cpu.f0.num\[31\] team_01_WB.instance_to_wrap.cpu.f0.num\[25\]
+ _04470_ _04585_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10387__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08044__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14117__A2 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08078_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] team_01_WB.instance_to_wrap.cpu.K0.keyvalid
+ _04523_ _04552_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout881_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10139__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12205__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[0\] net962 vssd1
+ vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09544__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 _02061_ vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[26\] vssd1 vssd1 vccd1 vccd1
+ net1637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[6\] vssd1 vssd1 vccd1 vccd1
+ net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[25\] vssd1 vssd1 vccd1 vccd1
+ net1659 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13628__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold54 net159 vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 _03519_ vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08919__A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold76 team_01_WB.instance_to_wrap.cpu.f0.write_data\[15\] vssd1 vssd1 vccd1 vccd1
+ net1692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 net131 vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold98 team_01_WB.instance_to_wrap.cpu.LCD0.lcd_rs vssd1 vssd1 vccd1 vccd1 net1714
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ net1963 net292 net472 vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__mux2_1
XANTENNA__09741__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11345__A team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18093__1587 vssd1 vssd1 vccd1 vccd1 _18093__1587/HI net1587 sky130_fd_sc_hd__conb_1
X_13730_ team_01_WB.instance_to_wrap.cpu.DM0.state\[0\] _04132_ _04133_ net1161 vssd1
+ vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__a22o_1
X_10942_ _06636_ _06671_ _06707_ net372 net549 net539 vssd1 vssd1 vccd1 vccd1 _07282_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11472__A1_N net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10311__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11064__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13661_ _03874_ _03875_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10873_ net528 _07212_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__nor2_1
X_15400_ net1274 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12612_ net3259 net303 net395 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16380_ clknet_leaf_77_wb_clk_i net1806 _00363_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_130_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13592_ net982 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _04035_ _04036_
+ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15331_ net1186 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12543_ net2286 net230 net405 vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08373__B team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18050_ net1550 vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__buf_2
XFILLER_0_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15262_ net1251 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__inv_2
X_12474_ net2380 net259 net411 vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17645__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17001_ clknet_leaf_9_wb_clk_i _02688_ _00984_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14213_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] vssd1 vssd1 vccd1
+ vccd1 _02274_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15487__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11425_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] _07736_ vssd1 vssd1 vccd1 vccd1
+ _07737_ sky130_fd_sc_hd__nand2_1
X_15193_ net1258 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__inv_2
XANTENNA__10378__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_7 _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14144_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[103\] _04244_ _04245_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[87\]
+ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__a22o_1
X_11356_ _04483_ _07684_ vssd1 vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__nor2_1
XANTENNA__09783__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13316__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[18\] net951
+ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__and3_1
X_14075_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[44\] _04246_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[108\]
+ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__a22o_1
XANTENNA__12115__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17795__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11287_ _06961_ _07622_ _07625_ _07626_ vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__or4_1
X_13026_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[60\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[68\]
+ net856 vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__mux2_1
X_17903_ net1423 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_94_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10238_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[9\] net780 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_89_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_0__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1030 net1031 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11954__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1041 net1045 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_23_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10169_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[10\] net790 net750 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__a22o_1
X_17834_ clknet_leaf_75_wb_clk_i net2543 _01774_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[104\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1052 net1053 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1063 team_01_WB.instance_to_wrap.cpu.f0.i\[22\] vssd1 vssd1 vccd1 vccd1 net1063
+ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08829__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1074 net1075 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1085 net1086 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__buf_1
XFILLER_0_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1096 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1
+ net1096 sky130_fd_sc_hd__buf_4
X_17765_ clknet_leaf_72_wb_clk_i net3167 _01705_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_14977_ net1246 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15950__A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13928_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__and2_2
XFILLER_0_72_1615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16716_ clknet_leaf_116_wb_clk_i _02403_ _00699_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_17696_ clknet_leaf_101_wb_clk_i _03380_ _01637_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10302__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16647_ clknet_leaf_16_wb_clk_i _02334_ _00630_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13859_ net1163 net1058 net3292 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[20\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_18_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13470__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16578_ clknet_leaf_32_wb_clk_i _02265_ _00561_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15529_ net1231 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09050_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[12\] net908
+ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10081__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09098__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08001_ net1067 vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold502 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10037__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold524 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09774__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold535 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09826__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold546 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold568 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09952_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[3\] net976 vssd1
+ vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11318__C1 _07650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08903_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[2\] net932 vssd1
+ vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__and3_1
XANTENNA__09526__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[5\] net963 vssd1
+ vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout295_A _07926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08734__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__A2 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2818 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[1\] net883 vssd1
+ vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__and3_1
Xhold1213 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2829 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1002_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1224 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[12\] vssd1 vssd1 vccd1 vccd1
+ net2840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1246 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2873 sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[4\] net680 _05078_ _05096_
+ net706 vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout462_A _07955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1268 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2895 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17518__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08696_ _05032_ _05033_ _05034_ _05035_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__or4_2
XFILLER_0_75_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10500__C net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10844__A1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12695__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1371_A net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout727_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17668__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08905__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09317_ net598 _05654_ _05656_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__o21a_2
XFILLER_0_36_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[21\] net675 net673 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10943__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09179_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[16\] net894 vssd1
+ vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11210_ _06903_ _07043_ _07548_ net554 vssd1 vssd1 vccd1 vccd1 _07550_ sky130_fd_sc_hd__a22o_1
X_12190_ _07790_ _07791_ net575 vssd1 vssd1 vccd1 vccd1 _07959_ sky130_fd_sc_hd__and3_4
XFILLER_0_47_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09736__C net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08640__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141_ net371 _07479_ _07480_ _07389_ vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__o31a_1
XFILLER_0_124_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11072_ _07403_ _07406_ _07407_ _07411_ _07364_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__a41o_1
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
XANTENNA__09517__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
X_10023_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[1\] net816 net805 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__a22o_1
X_14900_ net1312 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__inv_2
XANTENNA__11774__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15880_ net1382 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__inv_2
XANTENNA__10532__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14831_ net1214 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__inv_2
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09471__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17550_ clknet_leaf_6_wb_clk_i _03237_ _01533_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14762_ net1325 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11974_ net1892 net269 net471 vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16501_ clknet_leaf_108_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_read_i
+ _00484_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.READ_I sky130_fd_sc_hd__dfrtp_1
X_13713_ team_01_WB.instance_to_wrap.cpu.c0.count\[4\] _04101_ team_01_WB.instance_to_wrap.cpu.c0.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10925_ net527 _07215_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__nand2_1
X_17481_ clknet_leaf_10_wb_clk_i _03168_ _01464_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14693_ net1321 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16432_ clknet_leaf_104_wb_clk_i _02186_ _00415_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_141_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_141_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13644_ net723 _07323_ net1068 vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10856_ net337 net334 _07194_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__mux2_1
XANTENNA__08384__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16363_ clknet_leaf_86_wb_clk_i net2446 _00346_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13575_ net185 _04020_ _04021_ net725 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10787_ _04919_ net505 vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__xnor2_1
X_18102_ net1589 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15314_ net1235 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12526_ net2357 net216 net405 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__mux2_1
XANTENNA__11260__A1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16294_ clknet_leaf_68_wb_clk_i net2728 _00277_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18033_ net1533 vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__buf_2
XFILLER_0_124_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11949__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15245_ net1212 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__inv_2
X_12457_ net2118 net191 net413 vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15010__A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] _07700_ _07707_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\]
+ vssd1 vssd1 vccd1 vccd1 _07727_ sky130_fd_sc_hd__a31o_1
X_15176_ net1287 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__inv_2
X_17901__1421 vssd1 vssd1 vccd1 vccd1 _17901__1421/HI net1421 sky130_fd_sc_hd__conb_1
X_12388_ net2722 net316 net426 vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__mux2_1
XANTENNA__08550__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14127_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[30\] _04243_ _04254_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[102\]
+ _04412_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__a221o_1
X_11339_ _04469_ _04470_ vssd1 vssd1 vccd1 vccd1 _07668_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10771__B1 _07110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09943__A _05115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14058_ _04217_ _04260_ _04343_ _04346_ _04146_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__o41a_1
XFILLER_0_24_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11684__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[77\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[85\]
+ net855 vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__mux2_1
XANTENNA__13465__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17817_ clknet_leaf_77_wb_clk_i _03493_ _01757_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08550_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[19\] net897
+ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__and3_1
X_17748_ clknet_leaf_66_wb_clk_i _03424_ _01688_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16565__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10320__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10826__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08481_ net1004 net881 vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__and2_1
XANTENNA__17810__CLK clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08495__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09692__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17679_ clknet_leaf_94_wb_clk_i _03363_ _01620_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_134_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08294__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09102_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[13\] net906
+ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10054__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09995__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09033_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[9\] net705 _05370_ _05372_
+ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_87_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout210_A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout308_A _07935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09747__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold310 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold332 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold354 team_01_WB.instance_to_wrap.a1.ADR_I\[24\] vssd1 vssd1 vccd1 vccd1 net1970
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold365 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold376 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10762__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1217_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[47\] vssd1 vssd1 vccd1 vccd1
+ net2003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout801 _04646_ vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__buf_6
Xhold398 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09853__A _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09935_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[4\] net817 net755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__a22o_1
Xfanout812 net814 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__buf_4
Xfanout823 net824 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__buf_2
Xfanout834 team_01_WB.instance_to_wrap.cpu.RU0.next_ihit vssd1 vssd1 vccd1 vccd1 net834
+ sky130_fd_sc_hd__buf_2
XANTENNA_fanout677_A _04790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout845 net846 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__buf_2
XANTENNA__17340__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout856 net869 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__clkbuf_4
Xfanout867 net868 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__buf_2
X_09866_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[12\] net813 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10514__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout878 _04810_ vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_4
Xhold1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 net891 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__buf_4
XANTENNA__09380__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1032 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ net1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[1\] net937 vssd1
+ vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__and3_1
Xhold1043 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09291__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09797_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[14\] net953
+ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__and3_1
Xhold1054 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout844_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1065 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[11\] vssd1 vssd1 vccd1 vccd1
+ net2681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15590__A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2692 sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[4\] net909 vssd1
+ vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2714 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10230__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10817__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13822__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08679_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[7\] net901 vssd1
+ vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10710_ net529 _07049_ _06965_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11690_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[13\] _07553_ net717 vssd1 vssd1
+ vccd1 vccd1 _07889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08635__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11342__B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10641_ _06974_ _06977_ _06978_ net554 vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10045__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11242__A1 _05729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13360_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] net1064 vssd1 vssd1 vccd1 vccd1
+ _03831_ sky130_fd_sc_hd__xor2_1
XANTENNA__09986__A2 _04684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10572_ _04746_ _06910_ vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__or2_2
XANTENNA__08932__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12311_ net2235 net289 net433 vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__mux2_1
XANTENNA__11769__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13291_ net2396 net825 _03775_ _03777_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15030_ net1247 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__inv_2
X_12242_ net2810 net234 net441 vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12742__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ net1841 net263 net449 vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11124_ _07451_ _07459_ _07462_ _07463_ vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__nor4_1
X_16981_ clknet_leaf_125_wb_clk_i _02668_ _00964_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11055_ net557 _06280_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15932_ net1388 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__inv_2
XANTENNA__10505__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09371__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16588__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[1\] net809 _06345_ vssd1
+ vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__a21o_1
XANTENNA__09910__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15863_ net1385 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17602_ clknet_leaf_70_wb_clk_i _03289_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_14814_ net1274 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__inv_2
X_15794_ net1381 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10808__A1 _07015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17533_ clknet_leaf_49_wb_clk_i _03220_ _01516_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14745_ net1311 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_103_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11957_ net2171 _07941_ net476 vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10908_ _06984_ _07000_ net517 vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__mux2_1
X_17464_ clknet_leaf_25_wb_clk_i _03151_ _01447_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10284__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14676_ net1374 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ net2222 net305 net485 vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09003__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16415_ clknet_leaf_86_wb_clk_i _02169_ _00398_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13627_ net187 _04064_ _04065_ net728 vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__a211o_1
XANTENNA__11252__B _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10839_ _05491_ _06159_ _07177_ _07178_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17395_ clknet_leaf_135_wb_clk_i _03082_ _01378_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09426__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16346_ clknet_leaf_61_wb_clk_i _02100_ _00329_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[69\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_54_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09977__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13558_ net197 net193 _07815_ _07865_ net643 vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_137_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17213__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11679__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12509_ net2320 net287 net409 vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16277_ clknet_leaf_82_wb_clk_i _02031_ _00260_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13489_ _03949_ _03843_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_129_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18016_ net1516 vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_hd__buf_2
X_15228_ net1173 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11536__A2 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17363__CLK clknet_leaf_137_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15159_ net1200 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10315__C net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09673__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07981_ team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1 _04479_
+ sky130_fd_sc_hd__inv_2
XANTENNA__17890__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[21\] net819 net818 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12303__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09901__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[23\] net785 net775 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08602_ _04920_ _04940_ _04941_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09582_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[25\] net754 net745 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_121_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09114__A0 _05418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13997__B1 _04288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08533_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[18\] net660 _04853_
+ _04861_ _04864_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout258_A _07892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08464_ net1083 net881 vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__and2_1
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08455__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09417__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08395_ _04708_ _04716_ net714 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1
+ vccd1 vccd1 _04735_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout425_A _07966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09968__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08752__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1334_A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08471__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17706__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14174__B1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09016_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[9\] net927 vssd1
+ vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__and3_1
XANTENNA__09286__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout794_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11527__A2 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold140 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[0\] vssd1 vssd1 vccd1 vccd1
+ net1756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold151 net101 vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[10\] vssd1 vssd1 vccd1 vccd1
+ net1778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold173 team_01_WB.instance_to_wrap.cpu.f0.write_data\[20\] vssd1 vssd1 vccd1 vccd1
+ net1789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold184 _02023_ vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[2\] vssd1 vssd1 vccd1 vccd1 net1811
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16730__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13817__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout631 net635 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_4
X_09918_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[4\] net795 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__a22o_1
Xfanout642 _03572_ vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12213__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout653 _04819_ vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__buf_8
XANTENNA__10522__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout664 _04806_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_6
Xfanout675 _04791_ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__buf_6
XANTENNA__09353__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout686 _04780_ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__buf_4
XFILLER_0_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09849_ net377 _05378_ net561 vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__a21oi_1
Xfanout697 _04766_ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__buf_6
XANTENNA__11160__A0 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12860_ net2101 net296 net381 vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux2_1
XANTENNA__16880__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08927__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13988__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11811_ net1856 net288 net493 vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09656__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12791_ team_01_WB.instance_to_wrap.a1.ADR_I\[13\] net640 net607 _03622_ vssd1 vssd1
+ vccd1 vccd1 _02236_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17900__1420 vssd1 vssd1 vccd1 vccd1 _17900__1420/HI net1420 sky130_fd_sc_hd__conb_1
XFILLER_0_84_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14530_ net1394 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__inv_2
X_11742_ net1844 net309 net501 vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14461_ net1369 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__inv_2
X_11673_ _07812_ _07875_ vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__and2b_1
XFILLER_0_138_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13204__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16200_ clknet_leaf_114_wb_clk_i _01960_ _00188_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13412_ _04501_ _05224_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__or2_1
X_17180_ clknet_leaf_31_wb_clk_i _02867_ _01163_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09959__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ net554 _06858_ _06921_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__a21o_1
X_14392_ net1309 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16131_ clknet_leaf_93_wb_clk_i _00022_ _00119_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12963__B2 _03716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13343_ net585 _07688_ _03817_ net830 vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__a31o_1
XANTENNA__16260__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10555_ net545 net513 vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16062_ clknet_leaf_88_wb_clk_i _01855_ _00050_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_13274_ net1062 _03754_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__xnor2_1
X_10486_ _05870_ _05901_ _05869_ vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09196__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15013_ net1205 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12225_ _07794_ _07945_ net574 vssd1 vssd1 vccd1 vccd1 _07962_ sky130_fd_sc_hd__and3_4
XANTENNA__10726__A0 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08395__B2 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12156_ net2957 net292 net453 vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__mux2_1
XANTENNA__09924__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ _06905_ _07284_ _07446_ vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12123__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12087_ net2976 net305 net461 vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__mux2_1
X_16964_ clknet_leaf_54_wb_clk_i _02651_ _00947_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13140__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08147__B2 _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11038_ _07271_ _07272_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__nand2_1
X_15915_ net1402 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__inv_2
XANTENNA__08698__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16895_ clknet_leaf_26_wb_clk_i _02582_ _00878_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11962__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15846_ net1363 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13979__B1 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12989_ net2830 net1745 net867 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15777_ net1307 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17516_ clknet_leaf_132_wb_clk_i _03203_ _01499_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14728_ net1352 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14659_ net1381 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__inv_2
X_17447_ clknet_leaf_17_wb_clk_i _03134_ _01430_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16603__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08870__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10009__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09668__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08180_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[101\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[93\]
+ net1039 vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17378_ clknet_leaf_36_wb_clk_i _03065_ _01361_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13600__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12954__A1 _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11710__B net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16329_ clknet_leaf_64_wb_clk_i _02083_ _00312_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[52\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_116_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08622__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16753__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17879__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09583__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12033__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09703_ net1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[21\] net957
+ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__and3_1
XANTENNA__09335__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout375_A _06129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11872__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[23\] net962
+ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08747__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17259__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09565_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[25\] net963
+ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout542_A _05189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1284_A net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08466__B net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08516_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[18\] net926
+ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__and3_1
XANTENNA__11445__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09496_ _05808_ _05835_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08447_ net1087 net913 vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout807_A net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11323__D team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08378_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] _04711_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__or3b_1
XFILLER_0_74_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire328 _07574_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12945__A1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12208__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08613__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14147__B1 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10340_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[17\] net965
+ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10271_ net1120 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[19\] net943
+ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12010_ net2074 net259 net468 vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1404 net1414 vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__buf_2
Xfanout1415 net38 vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout450 _07958_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08129__A1 _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout461 _07955_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_50_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09326__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout472 _07952_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13961_ _04217_ _04220_ _04239_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_35_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout483 net484 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12878__S net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout494 _07944_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__buf_4
XFILLER_0_57_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11782__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15700_ net1293 vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__inv_2
X_12912_ net1619 net870 net357 _03683_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16680_ clknet_leaf_22_wb_clk_i _02367_ _00663_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09760__B net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13892_ _04139_ net571 _04197_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15631_ net1216 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__inv_2
X_12843_ net2753 net201 net379 vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__mux2_1
XANTENNA__10398__S net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16626__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10239__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15562_ net1278 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__inv_2
XANTENNA__11436__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12774_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] net1055 net364 _03610_
+ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14513_ net1398 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17301_ clknet_leaf_126_wb_clk_i _02988_ _01284_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11725_ net1915 net281 net501 vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__mux2_1
X_15493_ net1206 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17232_ clknet_leaf_126_wb_clk_i _02919_ _01215_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14444_ net1376 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11656_ net2824 net244 net499 vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16776__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08823__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12936__A1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11739__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10607_ net550 _06280_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17163_ clknet_leaf_5_wb_clk_i _02850_ _01146_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13594__D1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_86_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14375_ net1319 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12118__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08604__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11587_ _07803_ vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14138__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16114_ clknet_leaf_100_wb_clk_i _01889_ _00102_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13326_ _03798_ _03802_ _03804_ _00020_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__a2bb2o_1
X_17094_ clknet_leaf_42_wb_clk_i _02781_ _01077_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold909 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire884 _04803_ vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_2
X_10538_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[31\] net904
+ net659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[31\] vssd1 vssd1 vccd1
+ vccd1 _06878_ sky130_fd_sc_hd__a32o_1
XFILLER_0_126_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11957__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16045_ clknet_leaf_90_wb_clk_i net876 _00033_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.enable
+ sky130_fd_sc_hd__dfrtp_1
X_13257_ net1062 _03748_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__or2_1
XANTENNA__13738__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10469_ _06798_ _06800_ _06805_ _06808_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__or4_2
X_12208_ net2704 net261 net446 vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__mux2_1
X_13188_ net21 net835 net628 net1956 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12139_ net2228 net269 net454 vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__mux2_1
XANTENNA__10162__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17996_ net1496 vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__buf_2
XFILLER_0_104_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16156__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1609 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09951__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17401__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16947_ clknet_leaf_135_wb_clk_i _02634_ _00930_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13664__A2 _07489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16878_ clknet_leaf_6_wb_clk_i _02565_ _00861_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11705__B net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15829_ net1372 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17551__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09350_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[25\] net679 net654 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[25\]
+ _05686_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08301_ net1119 net966 vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_118_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09281_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[22\] net931 vssd1
+ vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08232_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[49\] net2023 net1053 vssd1 vssd1
+ vccd1 vccd1 _03455_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11440__B _07701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08163_ net2970 net2821 net1042 vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12028__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08094_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[17\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[16\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[19\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_77_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11867__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16024__A net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13352__A1 _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09564__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout492_A _07944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10072__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ _05324_ _05327_ net618 net617 vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__and4_1
XFILLER_0_122_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17081__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12698__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13655__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_A _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17914__1430 vssd1 vssd1 vccd1 vccd1 _17914__1430/HI net1430 sky130_fd_sc_hd__conb_1
XANTENNA__13383__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08477__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ _05935_ _05954_ _05955_ _05956_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__or4_1
XFILLER_0_74_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout924_A _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09548_ _05880_ _05885_ _05886_ _05887_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14080__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_120_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13830__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09479_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[30\] net683 _05817_
+ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_134_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08924__B net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11510_ net2429 net877 _07758_ _07782_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__o22a_1
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12490_ net3137 net189 net407 vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09739__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08643__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11441_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\] _07675_ net326 vssd1 vssd1 vccd1
+ vccd1 _07745_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08047__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14160_ _04195_ _04440_ net1411 vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13591__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11372_ net1065 _07676_ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__nand2_2
XFILLER_0_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08940__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11777__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13111_ net1 net844 vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__nor2_1
XANTENNA__10944__A3 _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10323_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[18\] net746 _06660_ _06661_
+ _06662_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_131_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14091_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[93\] _04240_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[125\]
+ _04377_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_128_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16179__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09547__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[44\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[52\]
+ net856 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__mux2_1
XANTENNA_input53_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_128_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10254_ net340 _06593_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09474__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1201 net1202 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__buf_4
Xfanout1212 net1214 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__buf_4
X_17850_ clknet_leaf_75_wb_clk_i net1996 _01790_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10185_ net582 _06521_ _06523_ _06524_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__a31o_4
Xfanout1223 net1227 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1234 net1235 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08770__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10413__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16801_ clknet_leaf_42_wb_clk_i _02488_ _00784_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1245 net1269 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__clkbuf_2
Xfanout1256 net1257 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__buf_4
X_17781_ clknet_leaf_72_wb_clk_i _03457_ _01721_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[51\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1267 net1268 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__buf_4
Xfanout1278 net1286 vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__buf_4
X_14993_ net1288 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__inv_2
Xfanout280 _07917_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_2
Xfanout291 net292 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__buf_2
Xfanout1289 net1294 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__buf_4
XANTENNA__17574__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16732_ clknet_leaf_32_wb_clk_i _02419_ _00715_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13944_ _04225_ _04234_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__nor2_4
XANTENNA__12401__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08818__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13875_ _04184_ _04185_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__a211o_1
X_16663_ clknet_leaf_136_wb_clk_i _02350_ _00646_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12826_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[2\] _07489_ net1034 vssd1 vssd1
+ vccd1 vccd1 _03647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11409__A1 _07701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15614_ net1263 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16594_ clknet_leaf_117_wb_clk_i _02281_ _00577_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14071__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12757_ net1970 net642 net606 _03599_ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__a22o_1
X_15545_ net1260 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10093__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11708_ net613 _07804_ _07903_ _07902_ vssd1 vssd1 vccd1 vccd1 _07904_ sky130_fd_sc_hd__a31o_4
XFILLER_0_72_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15476_ net1264 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12688_ net2163 net191 net385 vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09011__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14427_ net1366 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__inv_2
XANTENNA__08038__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17215_ clknet_leaf_7_wb_clk_i _02902_ _01198_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11639_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[24\] net715 net616 vssd1 vssd1
+ vccd1 vccd1 _07849_ sky130_fd_sc_hd__o21a_1
XANTENNA__10157__A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13582__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17146_ clknet_leaf_45_wb_clk_i _02833_ _01129_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09946__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14358_ net1363 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold706 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold717 team_01_WB.instance_to_wrap.a1.ADR_I\[28\] vssd1 vssd1 vccd1 vccd1 net2333
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold728 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ _07686_ _07709_ _03790_ net586 vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__o211a_1
X_17077_ clknet_leaf_124_wb_clk_i _02764_ _01060_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ net1385 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16028_ net1349 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__inv_2
X_08850_ _04755_ _05187_ _05188_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1406 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1417 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3033 sky130_fd_sc_hd__dlygate4sd3_1
X_08781_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[0\] net920 vssd1
+ vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__and3_1
X_17979_ net1479 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
Xhold1428 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1439 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3055 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13637__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11648__A1 _07154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11716__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08297__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16941__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09402_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[27\] net673 net668 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[27\]
+ _05738_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_62_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09069__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14062__A2 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08277__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09333_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[24\] net664 net659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10766__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout240_A _07870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_A _06911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10084__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09264_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[20\] net666 net653 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[20\]
+ _05603_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08215_ net2437 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[58\] net1043 vssd1 vssd1
+ vccd1 vccd1 _03472_ sky130_fd_sc_hd__mux2_1
XANTENNA__13558__D1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09195_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[17\] net919 vssd1
+ vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout505_A _06636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1247_A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09777__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ _04580_ _04581_ _04586_ _04587_ _04584_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17447__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09241__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08077_ _04515_ _04538_ _04544_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1414_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09294__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16471__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17597__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold11 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[6\] vssd1 vssd1 vccd1 vccd1 net1627
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold22 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[9\] vssd1 vssd1 vccd1 vccd1
+ net1638 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13825__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold33 team_01_WB.instance_to_wrap.cpu.f0.write_data\[29\] vssd1 vssd1 vccd1 vccd1
+ net1649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 net146 vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[8\] net690 _05316_ _05317_
+ _05318_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__a2111oi_1
Xhold55 net145 vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13628__A2 _07269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08919__B _05224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold66 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[1\] vssd1 vssd1 vccd1 vccd1
+ net1682 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12221__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold77 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[3\] vssd1 vssd1 vccd1 vccd1 net1693
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11990_ net2207 net317 net474 vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__mux2_1
Xhold88 _01996_ vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[5\] vssd1 vssd1 vccd1 vccd1 net1715
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08504__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08638__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11103__A3 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10941_ net526 _07280_ _07150_ _07062_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_97_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13660_ net982 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] _04091_ _04092_
+ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10872_ _07210_ _07211_ net518 vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__mux2_1
XANTENNA__08935__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12611_ net2538 net284 net398 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13591_ net723 _07611_ net1068 vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ net1313 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__inv_2
X_12542_ net1845 net287 net405 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09469__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09480__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15261_ net1252 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__inv_2
X_12473_ net2490 net233 net413 vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17000_ clknet_leaf_22_wb_clk_i _02687_ _00983_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14212_ net1760 vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13564__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ _04485_ _07701_ vssd1 vssd1 vccd1 vccd1 _07736_ sky130_fd_sc_hd__nor2_1
XANTENNA__09768__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15192_ net1172 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__inv_2
XANTENNA__09232__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14143_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[103\] _04254_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[111\]
+ _04427_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_39_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11355_ _04484_ _07683_ vssd1 vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16814__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10306_ _06642_ _06643_ _06644_ _06645_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__or4_1
X_14074_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[36\] _04230_ _04251_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[84\]
+ _04361_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11286_ _07019_ _07056_ _07111_ vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13025_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[61\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[69\]
+ net855 vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__mux2_1
X_17902_ net1422 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
X_10237_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[9\] net803 net751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_89_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1020 net1023 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_89_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1031 net1032 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09940__B1 _06278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1042 net1044 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_4
X_17833_ clknet_leaf_77_wb_clk_i net2828 _01773_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[103\]
+ sky130_fd_sc_hd__dfrtp_1
X_10168_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[10\] net819 _06506_
+ _06507_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1053 team_01_WB.instance_to_wrap.cpu.SR1.enable vssd1 vssd1 vccd1 vccd1 net1053
+ sky130_fd_sc_hd__buf_2
Xfanout1064 team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 net1064
+ sky130_fd_sc_hd__clkbuf_4
Xfanout1075 net1096 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_2
Xfanout1086 net1089 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__clkbuf_2
X_17764_ clknet_leaf_66_wb_clk_i _03440_ _01704_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12131__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1097 net1105 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__buf_4
X_10099_ _05264_ _05265_ _05301_ net378 vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__o31a_1
XFILLER_0_16_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14976_ net1244 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09006__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_63_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_117_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10838__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16715_ clknet_leaf_144_wb_clk_i _02402_ _00698_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08548__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13927_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__and2b_2
XFILLER_0_88_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13868__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17695_ clknet_leaf_99_wb_clk_i _03379_ _01636_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11970__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16646_ clknet_leaf_41_wb_clk_i _02333_ _00629_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13858_ net1163 net1058 net3285 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[19\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__14044__A2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12809_ net366 _03633_ _03634_ net1057 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__a32o_1
X_16577_ clknet_leaf_44_wb_clk_i _02264_ _00560_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13252__B1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13789_ _04154_ _04171_ _04172_ _04167_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a31o_1
XFILLER_0_130_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15528_ net1290 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15459_ net1188 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08000_ team_01_WB.instance_to_wrap.cpu.f0.num\[2\] vssd1 vssd1 vccd1 vccd1 _04498_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_4_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13555__A1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12814__B _07507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold503 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold514 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
X_17129_ clknet_leaf_8_wb_clk_i _02816_ _01112_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold525 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12306__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold536 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 net2152
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09951_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[3\] net955 vssd1
+ vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__and3_1
Xhold558 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold569 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[7\] vssd1 vssd1 vccd1 vccd1
+ net2185 sky130_fd_sc_hd__dlygate4sd3_1
X_08902_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[2\] net895 vssd1
+ vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09882_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[5\] net952 vssd1
+ vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09931__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08833_ net1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[1\] net911 vssd1
+ vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__and3_1
XANTENNA__08734__B2 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1203 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[97\] vssd1 vssd1 vccd1 vccd1
+ net2830 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10541__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1225 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2841 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1236 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2863 sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ _05100_ _05101_ _05102_ _05103_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__or4_1
XANTENNA__12041__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10350__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1258 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2874 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1269 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2885 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08458__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12294__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08695_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[7\] net658 _05014_ _05021_
+ _05024_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout455_A _07956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11880__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1197_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10844__A2 _07016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout622_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1364_A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10057__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09316_ net1111 net713 net600 net594 vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__a211o_1
XANTENNA__09998__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__C1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09289__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09247_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[21\] net700 _05586_ net706
+ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16837__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13546__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[16\] net691 _05515_ _05516_
+ _05517_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout991_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09214__A2 _04776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08129_ _04470_ team_01_WB.instance_to_wrap.cpu.f0.num\[25\] team_01_WB.instance_to_wrap.cpu.f0.num\[15\]
+ _04479_ _04598_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a221o_1
XANTENNA__12216__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11140_ net334 net338 _07390_ vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__mux2_1
XANTENNA__16987__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11071_ _07409_ _07410_ _07373_ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__a21bo_1
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__clkbuf_4
X_10022_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[1\] net742 _06359_ _06360_
+ _06361_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_60_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16217__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14830_ net1284 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14761_ net1329 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__inv_2
X_11973_ net1873 net236 net471 vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11790__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16500_ clknet_leaf_106_wb_clk_i _02254_ _00483_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10296__B1 _06634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10924_ net330 _07263_ _07262_ _07260_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13712_ net1632 _04504_ _03573_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__a21bo_1
X_17480_ clknet_leaf_30_wb_clk_i _03167_ _01463_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14692_ net1319 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14026__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17919__1607 vssd1 vssd1 vccd1 vccd1 net1607 _17919__1607/LO sky130_fd_sc_hd__conb_1
X_16431_ clknet_leaf_106_wb_clk_i _02185_ _00414_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10855_ net377 net331 vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__nor2_1
X_13643_ net187 _04077_ _04078_ net727 vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__a211o_1
XFILLER_0_116_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08384__B net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10048__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16362_ clknet_leaf_62_wb_clk_i _02116_ _00345_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[85\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13574_ net197 net193 _07876_ net643 vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__o211a_1
XANTENNA__09199__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10786_ _04919_ net505 net370 vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09453__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18101_ net638 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_1
X_15313_ net1324 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12525_ net3082 net222 net405 vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__mux2_1
X_16293_ clknet_leaf_76_wb_clk_i _02047_ _00276_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18032_ net1532 vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__buf_2
XFILLER_0_129_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12456_ _07790_ _07946_ net573 vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__and3_4
X_15244_ net1181 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_110_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08831__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ _07712_ _07726_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__nor2_1
X_15175_ net1328 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12387_ net2256 net318 net426 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__mux2_1
XANTENNA__12126__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14126_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[78\] _04235_ _04241_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[94\]
+ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__a22o_1
X_11338_ _07667_ net1756 _07655_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__mux2_1
XANTENNA__12760__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10771__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11965__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14057_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] _04237_ _04342_ _04344_
+ _04345_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__a2111o_1
X_11269_ _06903_ _06959_ vssd1 vssd1 vccd1 vccd1 _07609_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13008_ net2445 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[86\] net852 vssd1 vssd1
+ vccd1 vccd1 _02117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17142__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17816_ clknet_leaf_75_wb_clk_i net2590 _01756_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17747_ clknet_leaf_71_wb_clk_i _03423_ _01687_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14959_ net1212 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10287__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08480_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[23\] net893
+ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__and3_1
X_17678_ clknet_leaf_110_wb_clk_i net1159 _01619_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.pc_enable
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__14017__A2 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09692__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17888__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16629_ clknet_leaf_124_wb_clk_i _02316_ _00612_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08294__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11236__C1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09101_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[13\] net910
+ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__and3_1
X_09032_ _05363_ _05364_ _05365_ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__or4_2
XFILLER_0_32_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13528__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08741__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold300 net94 vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12036__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold311 team_01_WB.instance_to_wrap.cpu.f0.write_data\[11\] vssd1 vssd1 vccd1 vccd1
+ net1927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout203_A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold322 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10211__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold333 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[6\] vssd1 vssd1 vccd1 vccd1
+ net1960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold355 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 net1982
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11875__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net804 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold388 _03461_ vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[4\] net815 net739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold399 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[0\] vssd1 vssd1 vccd1 vccd1 net2015
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout813 net814 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__buf_6
Xfanout824 _04630_ vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__clkbuf_4
Xfanout835 _03737_ vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_4
Xfanout846 net848 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_2
Xfanout857 net859 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_4
X_09865_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[12\] net792 net789 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__a22o_1
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1000 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[58\] vssd1 vssd1 vccd1 vccd1
+ net2616 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09572__C net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout868 net869 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__buf_4
XANTENNA__11711__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 _04810_ vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__buf_2
Xhold1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08816_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[1\] net916 vssd1
+ vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__and3_1
Xhold1033 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10080__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09796_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[14\] net819 net753 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__a22o_1
Xhold1044 team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 net2660
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1055 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2693 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[4\] net888 vssd1
+ vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__and3_1
XANTENNA__17635__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1088 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1099 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[26\] vssd1 vssd1 vccd1 vccd1
+ net2715 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13391__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08678_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[7\] net907 vssd1
+ vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10817__A2 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14008__A2 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08485__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09683__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ net524 _06928_ vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09435__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11242__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10571_ _04746_ _06910_ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12310_ net2926 net255 net432 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__mux2_1
XANTENNA__13519__A1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13290_ net565 _03752_ _03776_ net829 vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08651__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12727__C1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12241_ net2495 net265 net440 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__mux2_1
XANTENNA__10255__A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12172_ net1906 net270 net447 vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__mux2_1
XANTENNA__11785__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ net516 _06957_ _07101_ vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__and3_1
XANTENNA__17165__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16980_ clknet_leaf_128_wb_clk_i _02667_ _00963_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11054_ _07062_ _07385_ _07391_ _07392_ _07393_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__a311o_1
X_15931_ net1402 vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10005_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[1\] net784 _04684_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15862_ net1385 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10421__C net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17601_ clknet_leaf_70_wb_clk_i _03288_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_14813_ net1262 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__inv_2
X_15793_ net1381 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__inv_2
X_17532_ clknet_leaf_31_wb_clk_i _03219_ _01515_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14744_ net1308 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__inv_2
X_11956_ net2911 net316 net478 vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08826__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10907_ net376 _06934_ _07014_ _07246_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__a31o_1
XANTENNA__13207__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17463_ clknet_leaf_140_wb_clk_i _03150_ _01446_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11887_ net2331 net312 net484 vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14675_ net1377 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16414_ clknet_leaf_79_wb_clk_i _02168_ _00397_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10838_ _05491_ net331 _07176_ _06912_ net369 vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__o221a_1
X_13626_ net199 net195 _07802_ _07907_ net645 vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_131_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17394_ clknet_leaf_134_wb_clk_i _03081_ _01377_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16345_ clknet_leaf_57_wb_clk_i _02099_ _00328_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[68\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10769_ net555 _07107_ _07108_ _06963_ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__o22a_1
X_13557_ _03925_ _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12508_ net2475 net258 net408 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
X_16276_ clknet_leaf_68_wb_clk_i _00004_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_4
X_13488_ _03844_ _03845_ _03946_ _05780_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__a32o_1
XFILLER_0_124_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10992__A1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18015_ net1515 vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_hd__buf_2
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08561__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12439_ net2597 net264 net417 vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__mux2_1
X_15227_ net1184 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09954__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15158_ net1202 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__inv_2
X_14109_ _04348_ _04395_ _04376_ net1169 vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15089_ net1292 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__inv_2
X_07980_ team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 _04478_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_59_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16532__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09650_ _05986_ _05987_ _05988_ _05989_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__or4_1
XFILLER_0_74_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08601_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[15\] net696 net652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09581_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[25\] net796 _05905_ _05907_
+ _05912_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_78_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09114__A1 _05453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16682__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08532_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[18\] net700 _04854_ _04860_
+ _04862_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_76_1390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08463_ net1106 net1109 net1115 net1113 vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_110_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08394_ net1156 _04717_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__nand2_1
XANTENNA__17038__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10059__B _06398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout320_A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08625__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_A _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10432__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09567__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09015_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[9\] net903 vssd1
+ vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10075__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1327_A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 _02144_ vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold141 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[27\] vssd1 vssd1 vccd1 vccd1
+ net1757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold152 _02002_ vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout787_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[22\] vssd1 vssd1 vccd1 vccd1
+ net1779 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__B2 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 team_01_WB.instance_to_wrap.a1.ADR_I\[29\] vssd1 vssd1 vccd1 vccd1 net1790
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13386__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17918__1606 vssd1 vssd1 vccd1 vccd1 net1606 _17918__1606/LO sky130_fd_sc_hd__conb_1
XFILLER_0_111_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold185 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[25\] vssd1 vssd1 vccd1 vccd1 net1801
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 _01968_ vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout610 _07685_ vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_2
Xfanout621 net622 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__buf_2
X_09917_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[4\] net788 net775 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[4\]
+ _06256_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__a221o_1
Xfanout632 net634 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout643 net644 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout954_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout654 _04819_ vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_4
Xfanout665 _04806_ vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout676 _04791_ vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__buf_4
X_09848_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] net627 _06186_ _06187_
+ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__a22o_2
Xfanout687 _04778_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__buf_6
XFILLER_0_77_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout698 _04763_ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__buf_8
XFILLER_0_38_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09779_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[15\] net796 net745 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11810_ net3110 net257 net493 vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15106__A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] net1056 net365 _03621_
+ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08646__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11741_ _07927_ _07928_ _07930_ net612 vssd1 vssd1 vccd1 vccd1 _07931_ sky130_fd_sc_hd__a22o_4
XANTENNA__11353__B team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_84_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14460_ net1348 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__inv_2
X_11672_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\]
+ _07809_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1 vccd1 vccd1
+ _07875_ sky130_fd_sc_hd__a31o_1
XANTENNA__08943__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09408__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10623_ net554 _06858_ _06921_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__a21oi_4
X_13411_ _03870_ _03871_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08616__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14391_ net1308 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_12__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_76_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_63_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10423__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13342_ _04481_ _07687_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__nand2_1
X_16130_ clknet_leaf_93_wb_clk_i _00021_ _00118_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12963__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10554_ _06890_ _06893_ net518 vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14165__A1 _04195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ _03749_ _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16061_ clknet_leaf_88_wb_clk_i _01854_ _00049_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_10485_ _06750_ _06819_ _06823_ _05902_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15012_ net1190 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__inv_2
XANTENNA__10416__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12224_ _07784_ _07789_ _07960_ vssd1 vssd1 vccd1 vccd1 _07961_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09041__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10726__A1 _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17800__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ net2106 net315 net453 vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__mux2_1
XANTENNA__12404__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11106_ net376 _07330_ _07445_ net531 vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__a22o_1
X_12086_ net3018 net310 net460 vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16963_ clknet_leaf_21_wb_clk_i _02650_ _00946_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13676__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11037_ _07375_ _07376_ _07374_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__a21oi_1
X_15914_ net1383 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__inv_2
XANTENNA__13140__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16894_ clknet_leaf_48_wb_clk_i _02581_ _00877_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09895__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15845_ net1363 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15776_ net1321 vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12988_ net2599 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[106\] net868 vssd1 vssd1
+ vccd1 vccd1 _02137_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09647__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09014__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08556__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17515_ clknet_leaf_4_wb_clk_i _03202_ _01498_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14727_ net1347 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__inv_2
X_11939_ net1947 net237 net475 vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14855__A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10662__A0 _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17446_ clknet_leaf_42_wb_clk_i _03133_ _01429_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09949__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14658_ net1381 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__inv_2
XANTENNA__08853__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08607__A0 _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13609_ net982 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _04049_ _04050_
+ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__a22o_1
X_17377_ clknet_leaf_43_wb_clk_i _03064_ _01360_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14589_ net1409 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16328_ clknet_leaf_73_wb_clk_i _02082_ _00311_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08083__A1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10965__A1 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16259_ clknet_leaf_104_wb_clk_i net1849 _00247_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10326__C net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17480__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12822__B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1053 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12314__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09702_ net1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[21\] net971
+ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__and3_1
XANTENNA__13131__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11142__A1 _05262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09633_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[23\] net945 vssd1
+ vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__and3_1
XANTENNA__12890__A1 _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout270_A _07877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09564_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[25\] net979
+ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_4_8__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14092__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08515_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[18\] net878
+ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_110_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_52_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09495_ _05833_ _05834_ net599 vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__mux2_2
XFILLER_0_81_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16428__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout535_A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1277_A net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08446_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[23\] net900
+ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13198__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08377_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] _04711_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout702_A _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12945__A2 _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16578__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09271__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09297__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09810__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17823__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15596__A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09594__A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ net1120 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[19\] net975
+ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__and3_1
XANTENNA__13828__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10708__A1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1405 net1413 vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__buf_4
XFILLER_0_100_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11348__B team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout440 _07962_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_4
XANTENNA__08003__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13122__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout451 net454 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_6
Xfanout462 _07955_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13960_ _04217_ _04220_ _04223_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_35_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout473 _07952_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_50_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11133__A1 _05189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout484 net486 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_6
XANTENNA__08938__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11133__B2 _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout495 net498 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_50_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12911_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[19\] _03682_ net1030 vssd1
+ vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13891_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__or2_1
XANTENNA__12881__A1 _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15630_ net1285 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12842_ net2889 net207 net379 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__mux2_1
XANTENNA__14083__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15561_ net1230 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__inv_2
XANTENNA__08837__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12773_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] _07251_ net1027 vssd1 vssd1
+ vccd1 vccd1 _03610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17300_ clknet_leaf_128_wb_clk_i _02987_ _01283_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ net1384 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _07913_ _07914_ _07916_ net613 vssd1 vssd1 vccd1 vccd1 _07917_ sky130_fd_sc_hd__a22o_4
X_15492_ net1239 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ clknet_leaf_143_wb_clk_i _02918_ _01214_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13189__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14443_ net1344 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__inv_2
X_11655_ net611 _07816_ _07861_ _07860_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__a31o_4
XFILLER_0_65_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10606_ net546 _06250_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__nor2_1
XANTENNA__12936__A2 _03699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17162_ clknet_leaf_2_wb_clk_i _02849_ _01145_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_88_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14374_ net1319 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__inv_2
X_11586_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\]
+ _07801_ vssd1 vssd1 vccd1 vccd1 _07803_ sky130_fd_sc_hd__and3_1
XANTENNA__09801__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16113_ clknet_leaf_99_wb_clk_i _01888_ _00101_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10537_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[31\] net663 net653 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[31\]
+ _06876_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__a221o_1
X_13325_ _07705_ _03803_ net828 vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17093_ clknet_leaf_38_wb_clk_i _02780_ _01076_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09000__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16044_ clknet_leaf_68_wb_clk_i _01838_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10468_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[26\] net796 net770 _06806_
+ _06807_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__a2111o_1
X_13256_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] _03747_ vssd1 vssd1 vccd1 vccd1
+ _03748_ sky130_fd_sc_hd__or2_1
XANTENNA__13738__B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12207_ net3021 net232 net445 vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__mux2_1
X_13187_ net22 net835 net628 net1697 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12134__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10399_ _05529_ _05730_ vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__xor2_1
XANTENNA__10175__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09009__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12138_ net2865 net235 net451 vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__mux2_1
X_17995_ net1495 vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10162__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09317__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11973__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08997__A1_N team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16946_ clknet_leaf_134_wb_clk_i _02633_ _00929_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12069_ net2884 net246 net459 vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08848__A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16877_ clknet_leaf_140_wb_clk_i _02564_ _00860_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12872__A1 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09670__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11274__A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15828_ net1373 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14074__B1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15759_ net1400 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__inv_2
XANTENNA__12624__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08300_ net1154 net1152 net1149 net1146 vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__and4b_1
XFILLER_0_115_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09280_ _05595_ _05619_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_118_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917__1605 vssd1 vssd1 vccd1 vccd1 net1605 _17917__1605/LO sky130_fd_sc_hd__conb_1
XANTENNA__08583__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08231_ net2481 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[42\] net1043 vssd1 vssd1
+ vccd1 vccd1 _03456_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17429_ clknet_leaf_124_wb_clk_i _03116_ _01412_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12309__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08162_ net2536 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[111\] net1046 vssd1 vssd1
+ vccd1 vccd1 _03525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08093_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[21\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[20\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[23\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13337__C1 _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08359__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12044__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10166__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17226__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[8\] net665 _05332_ _05333_
+ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__11883__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout485_A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11115__B2 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__A2 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12863__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1394_A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08477__B net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16250__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17376__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08531__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10874__A0 _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[24\] net741 _05937_ _05943_
+ _05948_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_92_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09547_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[28\] _04659_ net762
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[28\] vssd1 vssd1 vccd1 vccd1
+ _05887_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17929__1431 vssd1 vssd1 vccd1 vccd1 _17929__1431/HI net1431 sky130_fd_sc_hd__conb_1
XFILLER_0_4_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09478_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[30\] net665 net651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08924__C net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08429_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[23\] net922
+ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_43_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12219__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11440_ net327 _07701_ _07744_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08047__B2 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10929__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08598__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11371_ team_01_WB.instance_to_wrap.cpu.f0.i\[7\] team_01_WB.instance_to_wrap.cpu.f0.i\[6\]
+ _07675_ vssd1 vssd1 vccd1 vccd1 _07700_ sky130_fd_sc_hd__and3_2
XANTENNA__13591__A2 _07611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13110_ team_01_WB.instance_to_wrap.a1.curr_state\[2\] team_01_WB.instance_to_wrap.a1.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__or2_1
X_10322_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[18\] net969
+ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__and3_1
XANTENNA__13328__C1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14090_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[45\] _04256_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[109\]
+ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13041_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[45\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[53\]
+ net855 vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10253_ _05374_ _06592_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10184_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[10\] net767 vssd1 vssd1
+ vccd1 vccd1 _06524_ sky130_fd_sc_hd__nor2_1
XANTENNA_input46_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1202 net1203 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__clkbuf_4
Xfanout1213 net1214 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_33_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1224 net1227 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11793__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1235 net1236 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16800_ clknet_leaf_33_wb_clk_i _02487_ _00783_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08770__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1246 net1249 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__buf_4
X_17780_ clknet_leaf_66_wb_clk_i net2482 _01720_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17719__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11106__A1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14992_ net1272 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_135_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_135_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1257 net1261 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11106__B2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout270 _07877_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_2
Xfanout1268 net1269 vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__clkbuf_4
Xfanout1279 net1286 vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13500__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout281 _07917_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_2
X_16731_ clknet_leaf_50_wb_clk_i _02418_ _00714_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__buf_2
X_13943_ _04218_ _04234_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__nor2_4
XFILLER_0_96_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16662_ clknet_leaf_141_wb_clk_i _02349_ _00645_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13874_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1 _04185_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_9_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15613_ net1262 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
XANTENNA__16743__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ net2476 net640 net607 _03646_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a22o_1
X_16593_ clknet_leaf_123_wb_clk_i _02280_ _00576_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_69_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15544_ net1183 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__inv_2
X_12756_ net363 _03597_ _03598_ net1055 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__a32o_1
XANTENNA__08607__S _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08834__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\]
+ _07800_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1 vccd1 vccd1
+ _07903_ sky130_fd_sc_hd__a31o_1
X_15475_ net1278 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12129__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ _07791_ _07942_ net574 vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__and3_4
XFILLER_0_56_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17214_ clknet_leaf_44_wb_clk_i _02901_ _01197_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14426_ net1360 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09235__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11638_ net715 _07600_ vssd1 vssd1 vccd1 vccd1 _07848_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10157__B _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11968__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08589__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17145_ clknet_leaf_46_wb_clk_i _02832_ _01128_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14357_ net1364 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__inv_2
XANTENNA__13582__A2 _07541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11569_ net3170 net153 team_01_WB.instance_to_wrap.cpu.K0.next_state vssd1 vssd1
+ vccd1 vccd1 _03272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10396__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold707 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13319__C1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12790__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17249__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold718 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ net610 _07707_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1
+ vccd1 _03790_ sky130_fd_sc_hd__a21o_1
Xhold729 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[39\] vssd1 vssd1 vccd1 vccd1
+ net2345 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17076_ clknet_leaf_13_wb_clk_i _02763_ _01059_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14288_ net1368 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__inv_2
XANTENNA__09665__C net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16027_ net1362 vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__inv_2
XANTENNA__13334__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ net2603 net355 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1
+ vccd1 vccd1 _01911_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10148__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16273__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08761__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08780_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[0\] net660 _05117_ _05118_
+ _05119_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__a2111o_1
Xhold1407 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3023 sky130_fd_sc_hd__dlygate4sd3_1
X_17978_ net1478 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1418 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1429 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16929_ clknet_leaf_43_wb_clk_i _02616_ _00912_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17979__1479 vssd1 vssd1 vccd1 vccd1 _17979__1479/HI net1479 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_85_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08297__B net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10856__A0 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14047__B1 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09401_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[27\] net701 _04766_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10871__A3 _06065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09332_ _05665_ _05667_ _05669_ _05671_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__or4_1
XFILLER_0_87_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13270__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08744__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09263_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[20\] net692 net664 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12039__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout233_A net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10348__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08214_ net3097 net3064 net1051 vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09194_ net1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[17\] _04782_
+ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11878__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08145_ _04612_ _04613_ _04614_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout400_A _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10387__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1142_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12781__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08076_ _04525_ _04550_ _04551_ net569 net1929 vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__a32o_1
XANTENNA__13378__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10139__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1407_A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout867_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 _01972_ vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13394__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold23 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[4\] vssd1 vssd1 vccd1 vccd1
+ net1639 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12502__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08978_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[8\] net935 vssd1
+ vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__and3_1
Xhold34 team_01_WB.instance_to_wrap.a1.ADR_I\[5\] vssd1 vssd1 vccd1 vccd1 net1650
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 team_01_WB.instance_to_wrap.cpu.f0.write_data\[17\] vssd1 vssd1 vccd1 vccd1
+ net1661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 net1672
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16766__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[2\] vssd1 vssd1 vccd1 vccd1 net1683
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold78 _01969_ vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12836__A1 _07831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold89 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[26\] vssd1 vssd1 vccd1 vccd1
+ net1705 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08504__A2 _04837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10940_ _07059_ _07061_ net519 vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10311__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10942__S0 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10871_ net511 net510 _06032_ _06065_ net548 net537 vssd1 vssd1 vccd1 vccd1 _07211_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_45_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12610_ net2390 net252 net395 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__mux2_1
XANTENNA__08268__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13590_ net187 _04033_ _04034_ net728 vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_26_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08654__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11361__B team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_109_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12541_ net3046 net255 net403 vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15260_ net1171 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__inv_2
XANTENNA__16146__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12472_ net3117 net265 net411 vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11788__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14211_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\] vssd1 vssd1 vccd1
+ vccd1 _02276_ sky130_fd_sc_hd__clkbuf_1
X_11423_ _07701_ _07702_ _07735_ net326 vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15191_ net1196 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10378__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_9 _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14142_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[55\] _04236_ _04265_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11354_ net1064 net1065 vssd1 vssd1 vccd1 vccd1 _07683_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10705__B _05867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10305_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[18\] net819 net791 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08991__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14073_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[68\] _04233_ _04262_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[52\]
+ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__a22o_1
X_11285_ _07554_ _07566_ _07624_ vssd1 vssd1 vccd1 vccd1 _07625_ sky130_fd_sc_hd__or3_1
X_10236_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[9\] net786 net759 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[9\]
+ _06569_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13024_ net2359 net2262 net852 vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__mux2_1
X_17901_ net1421 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_0_30_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1010 net1013 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17916__1604 vssd1 vssd1 vccd1 vccd1 net1604 _17916__1604/LO sky130_fd_sc_hd__conb_1
Xfanout1021 net1022 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09940__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17832_ clknet_leaf_75_wb_clk_i _03508_ _01772_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[102\]
+ sky130_fd_sc_hd__dfrtp_1
X_10167_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[10\] net775 net772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__a22o_1
XANTENNA__12412__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1032 team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1 vccd1
+ net1032 sky130_fd_sc_hd__buf_2
Xfanout1043 net1044 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1054 net1055 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__buf_2
XFILLER_0_41_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1065 team_01_WB.instance_to_wrap.cpu.f0.i\[7\] vssd1 vssd1 vccd1 vccd1 net1065
+ sky130_fd_sc_hd__buf_2
XANTENNA__08829__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17763_ clknet_leaf_71_wb_clk_i _03439_ _01703_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[33\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1076 net1077 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__clkbuf_2
Xfanout1087 net1089 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__buf_2
XANTENNA__12827__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14975_ net1256 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__inv_2
X_10098_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] net626 _06436_ _06437_
+ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__a22o_4
Xfanout1098 net1100 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16714_ clknet_leaf_2_wb_clk_i _02401_ _00697_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13926_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__nand2b_4
XANTENNA__14029__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17694_ clknet_leaf_99_wb_clk_i _03378_ _01635_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_117_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10302__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16645_ clknet_leaf_31_wb_clk_i _02332_ _00628_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13857_ net1163 net1058 net3280 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[18\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_18_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12808_ net1033 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[7\] vssd1 vssd1 vccd1
+ vccd1 _03634_ sky130_fd_sc_hd__or2_1
X_16576_ clknet_leaf_30_wb_clk_i _02263_ _00559_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13252__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09456__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13788_ _04168_ _04170_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09022__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15527_ net1328 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_32_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12739_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] net1054 net363 _03586_
+ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__a22o_2
XFILLER_0_123_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09957__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15458_ net1312 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__inv_2
XANTENNA__08861__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17071__CLK clknet_leaf_143_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14409_ net1400 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13555__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13479__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15389_ net1250 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12763__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold504 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
X_17128_ clknet_leaf_24_wb_clk_i _02815_ _01111_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold515 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[13\] vssd1 vssd1 vccd1 vccd1 net2131
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold537 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[9\] vssd1 vssd1 vccd1 vccd1 net2164
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13307__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09950_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[3\] net950 vssd1
+ vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__and3_1
X_17059_ clknet_leaf_19_wb_clk_i _02746_ _01042_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold559 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08901_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[2\] net912 vssd1
+ vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09881_ _06165_ _06194_ _06220_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08832_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[1\] net911 vssd1
+ vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__and3_1
XANTENNA__12322__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10631__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1204 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1215 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2831 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10541__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1226 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2842 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1237 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2853 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08739__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1248 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2864 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[4\] net649 _05081_ _05085_
+ _05087_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__a2111o_1
Xhold1259 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[17\] vssd1 vssd1 vccd1 vccd1
+ net2875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08694_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[7\] net698 _05019_ _05022_
+ _05029_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_73_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1092_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout448_A _07958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09447__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17414__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10057__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08474__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09315_ net1111 net713 net594 vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10078__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1357_A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09246_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[21\] net682 net655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09177_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[16\] net885
+ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__and3_1
XANTENNA__13546__A2 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08128_ _04484_ team_01_WB.instance_to_wrap.cpu.f0.num\[9\] team_01_WB.instance_to_wrap.cpu.f0.num\[12\]
+ _04482_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_47_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout984_A _04499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08059_ _04514_ _04528_ _04529_ _04522_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_43_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11070_ _05006_ _06526_ _07374_ _06495_ _04969_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__o32a_1
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
X_10021_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[1\] net798 net792 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__a22o_1
XANTENNA__08725__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12232__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10532__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12809__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14760_ net1324 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__inv_2
XANTENNA__13482__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ net2553 net240 net471 vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__mux2_1
XANTENNA__09686__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08946__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13482__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18049__1549 vssd1 vssd1 vccd1 vccd1 _18049__1549/HI net1549 sky130_fd_sc_hd__conb_1
XANTENNA__09150__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ team_01_WB.instance_to_wrap.cpu.c0.count\[15\] _04502_ _04109_ _04125_ vssd1
+ vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[16\] sky130_fd_sc_hd__a31o_1
XANTENNA__10296__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10923_ _07212_ _07256_ net524 vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10687__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14691_ net1343 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16430_ clknet_leaf_96_wb_clk_i _02184_ _00413_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13642_ net200 net195 _07799_ _07920_ net645 vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_116_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10854_ net377 _06496_ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16361_ clknet_leaf_57_wb_clk_i _02115_ _00344_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[84\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_32_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13573_ _03918_ _04019_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10785_ net505 net335 net332 vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18100_ net637 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_1
X_15312_ net1224 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__inv_2
XANTENNA__10419__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12524_ net2253 net226 net403 vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ clknet_leaf_79_wb_clk_i _02046_ _00275_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08681__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18031_ net1531 vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__buf_2
X_15243_ net1298 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12455_ net2774 net293 net417 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__mux2_1
XANTENNA__09496__B _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12407__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17978__1478 vssd1 vssd1 vccd1 vccd1 _17978__1478/HI net1478 sky130_fd_sc_hd__conb_1
X_11406_ team_01_WB.instance_to_wrap.cpu.f0.i\[22\] _07694_ net325 vssd1 vssd1 vccd1
+ vccd1 _07726_ sky130_fd_sc_hd__o21ai_1
X_15174_ net1326 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__inv_2
X_12386_ net1962 net306 net426 vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__mux2_1
XANTENNA__16931__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14125_ _04405_ _04406_ _04408_ _04410_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__or4_1
X_11337_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] team_01_WB.instance_to_wrap.cpu.f0.state\[4\]
+ _04561_ _07652_ vssd1 vssd1 vccd1 vccd1 _07667_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14056_ _04226_ _04250_ _04255_ _04264_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__or4_1
X_11268_ _06915_ _07365_ _07366_ _06912_ _07607_ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__o221a_1
XANTENNA__13170__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13007_ net2435 net2327 net862 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__mux2_1
XANTENNA__12142__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10219_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[8\] net816 net769 _06557_
+ _06558_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11199_ net514 _07063_ _07099_ _07538_ vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09017__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17815_ clknet_leaf_61_wb_clk_i _03491_ _01755_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[85\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11981__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17746_ clknet_leaf_85_wb_clk_i _03422_ _01686_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14958_ net1282 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16311__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09141__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13909_ _04207_ net572 _04206_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__and3b_1
XFILLER_0_76_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10597__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17677_ clknet_leaf_111_wb_clk_i _03362_ _01618_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14889_ net1229 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11282__A _07088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16628_ clknet_leaf_12_wb_clk_i _02315_ _00611_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09429__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13225__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16559_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[25\]
+ _00542_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16461__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09100_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[13\] net899
+ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09031_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[9\] net700 _05348_ _05358_
+ net708 vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_60_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13528__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12317__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10626__A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11539__B2 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold301 _02025_ vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold312 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_29_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold323 team_01_WB.instance_to_wrap.cpu.f0.num\[0\] vssd1 vssd1 vccd1 vccd1 net1939
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 _03412_ vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold356 team_01_WB.instance_to_wrap.cpu.c0.count\[14\] vssd1 vssd1 vccd1 vccd1 net1972
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[23\] vssd1 vssd1 vccd1 vccd1
+ net1983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 team_01_WB.instance_to_wrap.cpu.c0.count\[2\] vssd1 vssd1 vccd1 vccd1 net1994
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[4\] net756 net750 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold389 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout803 net804 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_6
XFILLER_0_111_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout814 _04637_ vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__buf_4
Xfanout825 net828 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout398_A _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13161__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout836 _03737_ vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12052__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09864_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[12\] net803 net738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__a22o_1
Xfanout847 net848 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__buf_2
Xfanout858 net869 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__clkbuf_4
Xhold1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout869 _03718_ vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__buf_2
XANTENNA__10514__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1105_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11711__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[1\] net705 vssd1 vssd1
+ vccd1 vccd1 _05155_ sky130_fd_sc_hd__or2_1
XANTENNA__08469__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09380__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1023 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[21\] vssd1 vssd1 vccd1 vccd1 net2639
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _06134_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__inv_2
Xhold1034 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11891__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1045 _01914_ vssd1 vssd1 vccd1 vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1056 team_01_WB.instance_to_wrap.cpu.f0.num\[26\] vssd1 vssd1 vccd1 vccd1 net2672
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2683 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ net1008 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[4\] net888 vssd1
+ vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__and3_1
Xhold1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout732_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[7\] net900 vssd1
+ vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__and3_1
XANTENNA__10817__A3 _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08485__B net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11192__A _06598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_66_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_113_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17915__1603 vssd1 vssd1 vccd1 vccd1 net1603 _17915__1603/LO sky130_fd_sc_hd__conb_1
XFILLER_0_118_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09597__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10570_ _04736_ _04738_ vssd1 vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09840__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16954__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08932__C _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13519__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09229_ _04884_ _04919_ _05567_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__nor3_1
XANTENNA__12227__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12240_ net2276 net267 net439 vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10738__C1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12171_ net2301 net238 net447 vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08800__D1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11122_ net371 _07386_ _07388_ net338 _07461_ vssd1 vssd1 vccd1 vccd1 _07462_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold890 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13152__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11053_ _07388_ _06340_ net521 vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__and3b_1
X_15930_ net1331 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__inv_2
XANTENNA__10271__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10505__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16334__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[1\] net947 vssd1
+ vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09371__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15861_ net1396 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__inv_2
XANTENNA__11086__B net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17600_ clknet_leaf_70_wb_clk_i _03287_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_14812_ net1171 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__inv_2
X_15792_ net1317 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08676__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17531_ clknet_leaf_50_wb_clk_i _03218_ _01514_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1590 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[15\] vssd1 vssd1 vccd1 vccd1
+ net3206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14743_ net1308 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11955_ net3060 net320 net478 vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16484__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17462_ clknet_leaf_141_wb_clk_i _03149_ _01445_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10906_ _04884_ _06671_ _07244_ _07245_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_120_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08882__A1 _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13207__A1 net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14674_ net1377 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__inv_2
X_11886_ net2415 net296 net486 vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16413_ clknet_leaf_86_wb_clk_i _02167_ _00396_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_101_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11218__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13625_ _03892_ _04063_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__xnor2_1
X_10837_ net334 _07176_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__nand2_1
X_17393_ clknet_leaf_17_wb_clk_i _03080_ _01376_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09003__C _04799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09426__A3 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16344_ clknet_leaf_73_wb_clk_i net2092 _00327_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15302__A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13556_ _03923_ _03924_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__nor2_1
XANTENNA__09831__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768_ _06314_ _07055_ vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12507_ net3049 net261 net409 vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16275_ clknet_leaf_68_wb_clk_i _00003_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_124_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12137__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13487_ _03845_ _03946_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10699_ _06948_ _06953_ net534 vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18014_ net1514 vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_hd__buf_2
XFILLER_0_124_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15226_ net1189 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__inv_2
X_12438_ net2022 net268 net415 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11976__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15157_ net1222 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12369_ net3235 net272 net424 vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14108_ _04385_ _04394_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__or2_2
XFILLER_0_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09673__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15088_ net1270 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13143__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14039_ net1660 net605 _04328_ net1170 vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09362__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08600_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[15\] net689 _04923_
+ _04925_ _04926_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a2111o_1
XANTENNA__16827__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12600__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09580_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[25\] net787 net759 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[25\]
+ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08586__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08531_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[18\] net655 _04850_
+ _04855_ _04868_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13997__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17729_ clknet_leaf_100_wb_clk_i team_01_WB.instance_to_wrap.cpu.f0.next_write_i
+ _01669_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_i sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_100_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_54_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08462_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[23\] net922 vssd1
+ vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08393_ _04709_ _04732_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12957__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15212__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08752__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16207__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12047__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout313_A _07931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1055_A team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09014_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[9\] net924 vssd1
+ vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11886__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18048__1548 vssd1 vssd1 vccd1 vccd1 _18048__1548/HI net1548 sky130_fd_sc_hd__conb_1
XFILLER_0_79_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold120 team_01_WB.instance_to_wrap.cpu.f0.write_data\[18\] vssd1 vssd1 vccd1 vccd1
+ net1736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 team_01_WB.instance_to_wrap.cpu.f0.write_data\[24\] vssd1 vssd1 vccd1 vccd1
+ net1747 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1222_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold142 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[3\] vssd1 vssd1 vccd1 vccd1
+ net1758 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold153 net105 vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 _03436_ vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _02027_ vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout682_A _04787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold186 _01991_ vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 _04754_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10803__B net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout611 net614 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__buf_4
XANTENNA__13134__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09916_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[4\] net753 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout622 net624 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_4
Xfanout633 net634 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout644 _04839_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_4
Xfanout655 _04817_ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__buf_4
XANTENNA__10522__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout666 net667 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09353__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] net766 net623 vssd1
+ vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__o21a_1
Xfanout677 _04790_ vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__buf_6
XANTENNA__11696__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout688 _04776_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_6
Xfanout699 _04763_ vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12510__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13437__A1 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09778_ _06113_ _06114_ _06115_ _06117_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__or4_1
X_17977__1477 vssd1 vssd1 vccd1 vccd1 _17977__1477/HI net1477 sky130_fd_sc_hd__conb_1
XANTENNA__08927__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09105__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _05065_ _05066_ _05067_ _05068_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__or4_1
XANTENNA__13988__A2 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11740_ _07797_ _07929_ vssd1 vssd1 vccd1 vccd1 _07930_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10120__B1 _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11671_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[17\] _07232_ net716 vssd1 vssd1
+ vccd1 vccd1 _07874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15122__A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12948__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13410_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] _05220_ vssd1 vssd1 vccd1
+ vccd1 _03871_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10622_ _05839_ _06826_ _06828_ vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__nand3_1
XFILLER_0_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14390_ net1308 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09120__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13341_ _07681_ _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__nor2_1
X_10553_ _06891_ _06892_ net539 vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10266__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10974__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16060_ clknet_leaf_92_wb_clk_i _01853_ _00048_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_13272_ net1062 _03748_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10484_ _06750_ _06819_ _06823_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__a21o_1
XANTENNA__11796__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15011_ net1188 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12223_ _07790_ _07791_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] vssd1 vssd1
+ vccd1 vccd1 _07960_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12154_ net2183 net318 net452 vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__mux2_1
XANTENNA__08170__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13125__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ _07282_ _07285_ net516 vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16962_ clknet_leaf_35_wb_clk_i _02649_ _00945_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12085_ net2770 net296 net462 vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13676__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15913_ net1339 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__inv_2
X_11036_ _05006_ _06527_ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__or2_1
X_16893_ clknet_leaf_20_wb_clk_i _02580_ _00876_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15844_ net1351 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12420__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14201__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13979__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15775_ net1321 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__inv_2
X_12987_ net2496 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[107\] net865 vssd1 vssd1
+ vccd1 vccd1 _02138_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17514_ clknet_leaf_2_wb_clk_i _03201_ _01497_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14726_ net1352 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10111__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11938_ net2432 net242 net475 vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17445_ clknet_leaf_38_wb_clk_i _03132_ _01428_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10662__A1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14657_ net1237 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__inv_2
XANTENNA__10875__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11869_ net2315 net203 net483 vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12939__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13608_ net723 _07520_ net1068 vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__o21a_1
X_17376_ clknet_leaf_31_wb_clk_i _03063_ _01359_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14588_ net1393 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__inv_2
XANTENNA__09804__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13600__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09668__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16327_ clknet_leaf_67_wb_clk_i _02081_ _00310_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_116_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13539_ _03928_ _03931_ _03990_ _03927_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_116_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16258_ clknet_leaf_104_wb_clk_i net1622 _00246_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17625__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15209_ net1228 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10178__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16189_ clknet_leaf_115_wb_clk_i _01949_ _00177_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10904__A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09583__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13116__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17775__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10342__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ net1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[21\] net978
+ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__and3_1
XANTENNA__09335__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11142__A2 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[23\] net964
+ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__and3_1
XANTENNA__12330__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17005__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08747__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ net993 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[25\] net946 vssd1
+ vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__and3_1
XANTENNA__11454__B net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08514_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[18\] net915 vssd1
+ vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09494_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 net713 _04841_ vssd1 vssd1 vccd1
+ vccd1 _05834_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10653__A1 _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08445_ net1113 net1115 net1107 net1110 vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__and4bb_1
XANTENNA_fanout430_A _07965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17155__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1172_A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08376_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] _04715_ _04710_ vssd1 vssd1
+ vccd1 vccd1 _04716_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08482__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14781__A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14147__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout897_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13397__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12505__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10169__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1406 net1413 vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__buf_2
XFILLER_0_100_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13658__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11348__C net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout430 _07965_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout441 _07962_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_126_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09326__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout463 net464 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout474 _07952_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11133__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout485 net486 vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_50_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout496 net498 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12910_ _04918_ net578 net362 vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_31_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12240__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13890_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] net571 vssd1 vssd1 vccd1
+ vccd1 _03247_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_31_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12841_ net2524 net274 net380 vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__mux2_1
XANTENNA__10892__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15560_ net1287 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12772_ net1974 net641 net608 _03609_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__a22o_1
X_14511_ net1329 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _07800_ _07915_ vssd1 vssd1 vccd1 vccd1 _07916_ sky130_fd_sc_hd__nor2_1
X_15491_ net1189 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11380__A team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17230_ clknet_leaf_6_wb_clk_i _02917_ _01213_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14442_ net1376 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11654_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _07814_ vssd1 vssd1
+ vccd1 vccd1 _07861_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10605_ _06938_ _06944_ net518 vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__mux2_1
X_17161_ clknet_leaf_11_wb_clk_i _02848_ _01144_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14373_ net1349 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11585_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] _07801_ vssd1 vssd1 vccd1
+ vccd1 _07802_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16112_ clknet_leaf_90_wb_clk_i _01887_ _00100_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14138__A2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13324_ team_01_WB.instance_to_wrap.cpu.f0.i\[17\] _07703_ vssd1 vssd1 vccd1 vccd1
+ _03803_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_94_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17092_ clknet_leaf_52_wb_clk_i _02779_ _01075_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10536_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\] net665 net651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13346__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16043_ clknet_leaf_68_wb_clk_i _01837_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13255_ team_01_WB.instance_to_wrap.cpu.f0.i\[25\] team_01_WB.instance_to_wrap.cpu.f0.i\[24\]
+ _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__and3_1
X_10467_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[26\] net783 _06786_ _06788_
+ _06793_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12415__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12206_ net2796 net263 net443 vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_57_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13186_ net23 net835 net628 net1851 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__o22a_1
X_10398_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] _06737_ net622 vssd1
+ vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12137_ net2870 net240 net451 vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__mux2_1
X_17994_ net1494 vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__buf_2
XANTENNA__17028__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_109_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09317__A2 _05654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16945_ clknet_leaf_17_wb_clk_i _02632_ _00928_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12068_ net2966 net201 net459 vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__mux2_1
XANTENNA__09951__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08848__B _05153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12150__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15027__A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11019_ _07127_ _07358_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_105_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16876_ clknet_leaf_134_wb_clk_i _02563_ _00859_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08567__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15827_ net1373 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14866__A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18047__1547 vssd1 vssd1 vccd1 vccd1 _18047__1547/HI net1547 sky130_fd_sc_hd__conb_1
X_15758_ net1400 vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__inv_2
XANTENNA__08864__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14709_ net1305 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15689_ net1228 vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08230_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[51\] net3241 net1051 vssd1 vssd1
+ vccd1 vccd1 _03457_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17428_ clknet_leaf_11_wb_clk_i _03115_ _01411_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12388__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08161_ net1995 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[112\] net1052 vssd1 vssd1
+ vccd1 vccd1 _03526_ sky130_fd_sc_hd__mux2_1
XANTENNA__15697__A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17359_ clknet_leaf_0_wb_clk_i _03046_ _01342_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09695__A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08092_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid _04531_ vssd1 vssd1 vccd1 vccd1
+ _04563_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_77_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17976__1476 vssd1 vssd1 vccd1 vccd1 _17976__1476/HI net1476 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_77_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12325__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08994_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[8\] net896 vssd1
+ vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__and3_1
XANTENNA__10072__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1018_A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout380_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12060__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[24\] net748 _05938_ _05941_
+ _05944_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_39_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10874__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14776__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout645_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1387_A net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09546_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[28\] net805 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16545__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout812_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[30\] net673 net660 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08428_ net1084 net923 vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__and2_1
XANTENNA__08924__D net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13576__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09101__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[30\] net740 _04668_ _04664_
+ _04655_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_135_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11370_ net325 vssd1 vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08940__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10321_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[18\] net978 vssd1
+ vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__and3_1
XANTENNA__12235__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13040_ net2465 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[54\] net852 vssd1 vssd1
+ vccd1 vccd1 _02085_ sky130_fd_sc_hd__mux2_1
XANTENNA__09547__A2 _04659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10252_ net561 _05338_ _06564_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_128_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10183_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[10\] net753 _06522_
+ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__a21oi_1
Xfanout1203 net1204 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__clkbuf_2
Xfanout1214 net1218 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__buf_4
Xfanout1225 net1227 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__buf_4
Xfanout1236 net1415 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__clkbuf_4
X_14991_ net1216 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1247 net1249 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__buf_4
XANTENNA_input39_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout260 net261 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1258 net1261 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__buf_4
XANTENNA__16075__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout271 net272 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_2
XANTENNA__08507__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1269 net1415 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__clkbuf_4
Xfanout282 _07917_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_2
X_16730_ clknet_leaf_60_wb_clk_i _02417_ _00713_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13942_ _04222_ _04228_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__nand2_2
XANTENNA__17320__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout293 _07941_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__buf_2
XFILLER_0_92_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10865__A1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16661_ clknet_leaf_130_wb_clk_i _02348_ _00644_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13873_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__or4_1
XANTENNA__14686__A net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15612_ net1176 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
X_12824_ net365 _03644_ _03645_ net1057 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__a32o_1
X_16592_ clknet_leaf_122_wb_clk_i _02279_ _00575_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_74_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_104_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13264__C1 _04466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08684__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15543_ net1200 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12755_ net1027 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[24\] vssd1 vssd1 vccd1
+ vccd1 _03598_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ net720 _07531_ net615 _07901_ vssd1 vssd1 vccd1 vccd1 _07902_ sky130_fd_sc_hd__o211a_1
XANTENNA__10093__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15474_ net1233 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__inv_2
X_12686_ net2701 net292 net390 vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17213_ clknet_leaf_40_wb_clk_i _02900_ _01196_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14425_ net1374 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__inv_2
X_11637_ net2174 net210 net502 vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__mux2_1
XANTENNA__08038__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09011__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10157__C net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17144_ clknet_leaf_28_wb_clk_i _02831_ _01127_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14356_ net1375 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__inv_2
X_11568_ team_01_WB.instance_to_wrap.cpu.K0.count\[1\] team_01_WB.instance_to_wrap.cpu.K0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__nand2b_1
XANTENNA__09946__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold708 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13307_ net3238 net825 _03787_ _03789_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__o22a_1
XANTENNA__12790__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17075_ clknet_leaf_135_wb_clk_i _02762_ _01058_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10519_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[31\] net696 net662 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__a22o_1
Xhold719 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
X_14287_ net1374 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__inv_2
XANTENNA__12145__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11499_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[13\] _07756_ vssd1 vssd1 vccd1
+ vccd1 _07777_ sky130_fd_sc_hd__and2_1
X_16026_ net1363 vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__inv_2
X_13238_ net2919 net355 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1
+ vccd1 vccd1 _01912_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11984__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13765__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13169_ net137 net847 net842 net1803 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08859__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17977_ net1477 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_97_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1408 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1419 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16928_ clknet_leaf_33_wb_clk_i _02615_ _00911_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10305__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10856__A1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09710__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16859_ clknet_leaf_52_wb_clk_i _02546_ _00842_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09400_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[27\] net681 net659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_62_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09331_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[24\] net693 net649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[24\]
+ _05670_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10629__A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[20\] net695 _05600_
+ _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11281__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10084__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08213_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[68\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[60\]
+ net1041 vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09226__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09193_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[17\] net922 vssd1
+ vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout226_A _07827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08144_ team_01_WB.instance_to_wrap.cpu.f0.i\[30\] _04493_ _04496_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\]
+ _04590_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09777__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12781__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12055__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08075_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] _04524_ vssd1 vssd1 vccd1 vccd1
+ _04551_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1135_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap961 _04650_ vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_2
Xmax_cap972 _04635_ vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13097__D net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11894__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1302_A net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[81\] vssd1 vssd1 vccd1 vccd1 net1629
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[8\] net901 vssd1
+ vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__and3_1
Xhold24 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[5\] vssd1 vssd1 vccd1 vccd1
+ net1640 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout762_A _04674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 _02003_ vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 team_01_WB.instance_to_wrap.cpu.f0.write_data\[27\] vssd1 vssd1 vccd1 vccd1
+ net1662 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11195__A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold57 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[38\] vssd1 vssd1 vccd1 vccd1 net1673
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[14\] vssd1 vssd1 vccd1 vccd1
+ net1684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1
+ net1695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10870_ net507 _06636_ _06671_ _06707_ net548 net539 vssd1 vssd1 vccd1 vccd1 _07210_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08935__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09529_ net513 _05868_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09465__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12540_ net2578 net259 net404 vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10258__B _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08009__A team_01_WB.instance_to_wrap.cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_108_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12471_ net2571 net269 net413 vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14210_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] vssd1 vssd1 vccd1
+ vccd1 _02277_ sky130_fd_sc_hd__clkbuf_1
X_11422_ team_01_WB.instance_to_wrap.cpu.f0.i\[15\] _07689_ vssd1 vssd1 vccd1 vccd1
+ _07735_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_91_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15190_ net1201 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__inv_2
XANTENNA__09768__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08670__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14141_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[39\] _04230_ _04259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[23\]
+ _04425_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12772__B2 _03609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11353_ team_01_WB.instance_to_wrap.cpu.f0.i\[14\] team_01_WB.instance_to_wrap.cpu.f0.i\[13\]
+ _07679_ vssd1 vssd1 vccd1 vccd1 _07682_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10274__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10304_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[18\] net756 net735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14072_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[60\] _04258_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[20\]
+ _04359_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11284_ _07135_ _07611_ _07621_ _07623_ vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__or4_1
X_18046__1546 vssd1 vssd1 vccd1 vccd1 _18046__1546/HI net1546 sky130_fd_sc_hd__conb_1
XFILLER_0_24_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13023_ net2619 net2498 net861 vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__mux2_1
X_17900_ net1420 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
X_10235_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[9\] net818 _06573_ _06574_
+ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_89_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1000 net1001 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__buf_2
Xfanout1011 net1012 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17831_ clknet_leaf_62_wb_clk_i _03507_ _01771_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[101\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout1022 net1023 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_2
X_10166_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[10\] net747 net744 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__a22o_1
XANTENNA__09940__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1033 net1034 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__buf_2
Xfanout1044 net1045 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1055 team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1 vccd1
+ net1055 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1066 net1067 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__clkbuf_4
X_17762_ clknet_leaf_76_wb_clk_i net2457 _01702_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[32\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1077 net1078 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__clkbuf_2
Xfanout1088 net1089 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__buf_1
X_14974_ net1251 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__inv_2
X_10097_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] net765 net622 vssd1
+ vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__o21a_1
Xfanout1099 net1100 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__buf_1
XFILLER_0_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16713_ clknet_leaf_8_wb_clk_i _02400_ _00696_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13925_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__and2b_2
XANTENNA__14029__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10838__B2 _06912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09006__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17693_ clknet_leaf_99_wb_clk_i _03377_ _01634_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12929__A team_01_WB.instance_to_wrap.cpu.f0.write_data\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16644_ clknet_leaf_17_wb_clk_i _02331_ _00627_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13856_ net1163 net1058 net2080 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[17\]
+ sky130_fd_sc_hd__and3b_1
X_17975__1475 vssd1 vssd1 vccd1 vccd1 _17975__1475/HI net1475 sky130_fd_sc_hd__conb_1
XFILLER_0_92_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09303__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12807_ net1033 _07308_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13787_ _04168_ _04170_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__or2_1
X_16575_ clknet_leaf_24_wb_clk_i _02262_ _00558_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_130_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10999_ _07062_ _07338_ _07337_ _07333_ vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15526_ net1326 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__inv_2
X_12738_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[29\] _07056_ net1025 vssd1 vssd1
+ vccd1 vccd1 _03586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11979__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15457_ net1243 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__inv_2
X_12669_ net2062 net267 net387 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14408_ net1332 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_72_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15388_ net1174 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12763__B2 _03603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14339_ net1377 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__inv_2
X_17127_ clknet_leaf_15_wb_clk_i _02814_ _01110_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold505 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17366__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold516 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold527 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold538 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
X_17058_ clknet_leaf_35_wb_clk_i _02745_ _01041_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold549 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12515__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08900_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[2\] net937 vssd1
+ vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16009_ net1385 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__inv_2
X_09880_ _06218_ _06219_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__nand2_1
XANTENNA__12603__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10526__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09392__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16390__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08831_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[1\] net894 vssd1
+ vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__and3_1
XANTENNA__09931__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1205 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[110\] vssd1 vssd1 vccd1 vccd1
+ net2821 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10631__B net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1216 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2843 sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[4\] net675 _05086_ _05093_
+ _05099_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__a2111o_1
Xhold1238 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2865 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10350__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10829__A1 _07064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08693_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[7\] net679 _05010_ _05017_
+ _05028_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_135_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11743__A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08755__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1085_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] net702 _05648_ _05653_
+ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__o22a_4
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10057__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09998__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__B2 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11889__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09245_ _05578_ _05580_ _05584_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__or3_1
XANTENNA_hold1193_A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout510_A _05996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08771__B net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1252_A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09176_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[16\] net914 vssd1
+ vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08127_ _04468_ team_01_WB.instance_to_wrap.cpu.f0.num\[27\] team_01_WB.instance_to_wrap.cpu.f0.num\[24\]
+ _04471_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10765__A0 _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09883__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08058_ net1862 net569 _04525_ _04535_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12513__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__B1 _06855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10020_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[1\] net754 net749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__a22o_1
XANTENNA__09383__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13852__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ net1744 net273 net473 vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_95_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08489__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10915__S1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13710_ team_01_WB.instance_to_wrap.cpu.c0.count\[16\] _04111_ _04119_ vssd1 vssd1
+ vccd1 vccd1 _04125_ sky130_fd_sc_hd__and3_1
X_10922_ _06904_ _07261_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__nor2_1
XANTENNA__10296__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14690_ net1344 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13641_ _03865_ _03881_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__xnor2_1
X_10853_ _06530_ _07191_ _06501_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10269__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16360_ clknet_leaf_74_wb_clk_i _02114_ _00343_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10048__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13572_ _03857_ _03858_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__and2b_1
XANTENNA__08962__A _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10784_ _06893_ _06938_ net517 vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15311_ net1215 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11799__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12523_ net2428 net191 net403 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
X_16291_ clknet_leaf_86_wb_clk_i net1718 _00274_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16263__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17389__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18030_ net1530 vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__buf_2
X_15242_ net1277 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12454_ net2671 net314 net418 vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12745__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11405_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] _07712_ _07713_ net325 vssd1 vssd1
+ vccd1 vccd1 _03386_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15173_ net1208 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12385_ net2835 net310 net425 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14124_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[38\] _04221_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[118\]
+ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__a221o_1
XANTENNA__09793__A _06129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11336_ _07666_ net1809 _07655_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14055_ _04230_ _04243_ _04249_ _04256_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__or4_1
X_11267_ _04948_ _07606_ vssd1 vssd1 vccd1 vccd1 _07607_ sky130_fd_sc_hd__nand2_1
XANTENNA__10508__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13006_ net1633 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[88\] net860 vssd1 vssd1
+ vccd1 vccd1 _02119_ sky130_fd_sc_hd__mux2_1
XANTENNA__09374__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10218_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[8\] net757 _06539_ _06540_
+ _06546_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11547__B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11198_ _07100_ _07280_ _07361_ _07537_ _07535_ vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__a221o_1
XANTENNA__11181__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17814_ clknet_leaf_56_wb_clk_i _03490_ _01754_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[84\]
+ sky130_fd_sc_hd__dfstp_1
X_10149_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[11\] net755 net732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17745_ clknet_leaf_79_wb_clk_i net3207 _01685_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14957_ net1207 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13908_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\]
+ _04204_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__and3_1
XANTENNA__10287__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17676_ clknet_leaf_111_wb_clk_i _03361_ _01617_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14888_ net1274 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
XANTENNA__08575__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11282__B _07154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10692__C1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16627_ clknet_leaf_129_wb_clk_i _02314_ _00610_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13839_ net1165 net1061 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[0\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[0\] sky130_fd_sc_hd__and3b_1
XFILLER_0_130_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16606__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11236__B2 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16558_ clknet_leaf_115_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[24\]
+ _00541_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15509_ net1225 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16489_ clknet_leaf_103_wb_clk_i _02243_ _00472_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09030_ _05366_ _05367_ _05368_ _05369_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__or4_1
XFILLER_0_115_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16756__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12736__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold302 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[21\] vssd1 vssd1 vccd1 vccd1
+ net1918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 team_01_WB.instance_to_wrap.cpu.f0.write_data\[4\] vssd1 vssd1 vccd1 vccd1
+ net1929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10345__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10211__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold324 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[126\] vssd1 vssd1 vccd1 vccd1
+ net1940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold335 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold357 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ _06268_ _06269_ _06270_ _06271_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__or4_1
Xhold368 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 net1984
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[120\] vssd1 vssd1 vccd1 vccd1
+ net1995 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12333__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout804 _04643_ vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout815 net816 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__buf_6
XANTENNA__09365__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout826 net827 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09208__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09904__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09863_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[12\] net822 net762 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__a22o_1
Xfanout837 _03736_ vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__clkbuf_4
Xfanout848 _03731_ vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11172__B1 _06912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout293_A _07941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net869 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__clkbuf_2
Xhold1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
X_08814_ _04708_ net729 net720 _04838_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__o41a_2
XANTENNA__11711__A2 _07269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ _06129_ _06131_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1000_A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1035 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10080__C net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1046 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08745_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[4\] net925 vssd1
+ vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__and3_1
Xhold1057 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2684 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout460_A _07955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08258__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[7\] net919 vssd1
+ vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11192__B _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16286__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout725_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18045__1545 vssd1 vssd1 vccd1 vccd1 _18045__1545/HI net1545 sky130_fd_sc_hd__conb_1
XANTENNA__17531__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13621__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1575_A team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12508__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09228_ _04970_ _05379_ _05494_ _05567_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__nor4_2
XFILLER_0_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17681__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09159_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[16\] net648 _05496_
+ _05497_ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_115_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12170_ net1867 net241 net447 vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13847__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17974__1474 vssd1 vssd1 vccd1 vccd1 _17974__1474/HI net1474 sky130_fd_sc_hd__conb_1
XFILLER_0_62_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11121_ net526 _07460_ vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__nor2_1
XANTENNA__12243__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold880 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[99\] vssd1 vssd1 vccd1 vccd1
+ net2496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold891 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09118__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11052_ net526 _06313_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10003_ _06340_ _06342_ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__nor2_1
X_15860_ net1385 vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__inv_2
XANTENNA__14101__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17061__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14811_ net1184 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__inv_2
X_15791_ net1318 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__inv_2
Xhold1580 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3196 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11383__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17530_ clknet_leaf_60_wb_clk_i _03217_ _01513_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11954_ net2489 net308 net478 vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__mux2_1
Xhold1591 _03421_ vssd1 vssd1 vccd1 vccd1 net3207 sky130_fd_sc_hd__dlygate4sd3_1
X_14742_ net1308 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__inv_2
XANTENNA__08168__S net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10905_ _04884_ net332 _07243_ net335 net370 vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__a221o_1
X_14673_ net1382 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__inv_2
X_17461_ clknet_leaf_124_wb_clk_i _03148_ _01444_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11885_ net2968 net300 net485 vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13207__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08882__A2 _05219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11218__A1 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13624_ _03893_ _04051_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__nand2b_1
X_16412_ clknet_leaf_95_wb_clk_i _02166_ _00395_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10836_ _05491_ _06159_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_101_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17392_ clknet_leaf_15_wb_clk_i _03079_ _01375_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16779__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16343_ clknet_leaf_67_wb_clk_i net2193 _00326_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[66\]
+ sky130_fd_sc_hd__dfrtp_1
X_13555_ net980 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _04004_ _04005_
+ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__a22o_1
XANTENNA__12418__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10977__A0 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10767_ net524 _07106_ _06965_ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11322__S _07655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12506_ net2888 net232 net409 vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__mux2_1
X_16274_ clknet_leaf_67_wb_clk_i _00002_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_13486_ _03846_ _03847_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ _07036_ _07037_ net520 vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18013_ net1513 vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_hd__buf_2
X_15225_ net1259 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12437_ net2147 net237 net415 vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09595__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15156_ net1291 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12368_ net3219 net244 net423 vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09954__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14107_ _04387_ _04389_ _04391_ _04393_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11319_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] net1162 vssd1 vssd1 vccd1
+ vccd1 _07656_ sky130_fd_sc_hd__and2_1
X_15087_ net1215 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__inv_2
XANTENNA__12153__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12299_ net1934 net274 net433 vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__mux2_1
XANTENNA__13143__A1 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09347__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14038_ _04319_ _04325_ _04326_ _04327_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__or4_2
XANTENNA__17404__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08867__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15989_ net1407 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17554__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08530_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[18\] net889
+ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__and3_1
X_17728_ clknet_leaf_66_wb_clk_i _03405_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08461_ net1011 net923 vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17659_ clknet_leaf_90_wb_clk_i _03344_ _01600_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08873__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09698__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08392_ net1155 _04713_ net710 vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12957__B2 _03713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08625__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12328__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10432__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09013_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[9\] net937 vssd1
+ vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout306_A _07935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1048_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10075__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09586__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 _02012_ vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold121 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1
+ net1737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold132 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[7\] vssd1 vssd1 vccd1 vccd1
+ net1748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold143 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[19\] vssd1 vssd1 vccd1 vccd1
+ net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _02006_ vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12063__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold165 team_01_WB.instance_to_wrap.cpu.f0.write_data\[25\] vssd1 vssd1 vccd1 vccd1
+ net1781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 team_01_WB.instance_to_wrap.a1.ADR_I\[11\] vssd1 vssd1 vccd1 vccd1 net1792
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1215_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout601 _04754_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_4
Xhold187 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[7\] vssd1 vssd1 vccd1 vccd1 net1803
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 team_01_WB.instance_to_wrap.cpu.f0.write_data\[3\] vssd1 vssd1 vccd1 vccd1
+ net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 net614 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_4
X_09915_ _06250_ _06253_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__or2_2
XFILLER_0_10_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout623 net624 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout634 net635 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__buf_2
XANTENNA_fanout675_A _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 net646 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_4
Xfanout656 _04817_ vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_8
X_09846_ _06178_ _06185_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__or2_2
Xfanout667 _04804_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__buf_6
XANTENNA__11696__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08777__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout678 _04790_ vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__clkbuf_4
Xfanout689 _04773_ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_8
X_09777_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[15\] net813 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[15\]
+ _06116_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_124_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13437__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08728_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[5\] net695 _05046_ _05053_
+ _05059_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_96_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16921__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10656__C1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08659_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[10\] net691 _04986_ _04988_
+ _04991_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_96_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11670_ net1942 net236 net499 vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12948__A1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08943__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10621_ _06886_ _06887_ _06960_ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_137_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08616__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12238__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13340_ team_01_WB.instance_to_wrap.cpu.f0.i\[13\] _07679_ net566 vssd1 vssd1 vccd1
+ vccd1 _03815_ sky130_fd_sc_hd__o21ai_1
X_10552_ net505 _06671_ net544 vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__mux2_1
XANTENNA__10423__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13271_ net1652 _03761_ net825 vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10483_ _06781_ _06815_ _06822_ _06818_ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_129_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15010_ net1312 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__inv_2
X_12222_ net3124 net292 net444 vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__mux2_1
XANTENNA__09577__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13373__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_input69_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17427__CLK clknet_leaf_137_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09041__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12153_ net2042 net306 net452 vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11104_ _07064_ net329 _07395_ _07443_ vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__a22oi_1
XANTENNA__09329__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12084_ net2278 net299 net462 vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__mux2_1
X_16961_ clknet_leaf_48_wb_clk_i _02648_ _00944_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13676__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15912_ net1336 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__inv_2
X_11035_ _05006_ _06527_ vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12701__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16892_ clknet_leaf_39_wb_clk_i _02579_ _00875_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15843_ net1351 vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__inv_2
XANTENNA__11825__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12986_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[100\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[108\]
+ net858 vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__mux2_1
X_15774_ net1320 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17513_ clknet_leaf_9_wb_clk_i _03200_ _01496_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ net1346 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09014__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11937_ net2084 _07866_ net477 vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_45 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12937__A _04968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15313__A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17444_ clknet_leaf_53_wb_clk_i _03131_ _01427_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14656_ net1186 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__inv_2
X_11868_ net1788 net208 net483 vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09949__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08853__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10819_ net530 _07158_ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__nor2_1
XANTENNA__12939__B2 _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13607_ net187 _04047_ _04048_ net728 vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__a211o_1
XANTENNA__12148__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17375_ clknet_leaf_8_wb_clk_i _03062_ _01358_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14587_ net1408 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11799_ net2979 net276 net492 vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__mux2_1
XANTENNA__13600__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16326_ clknet_leaf_68_wb_clk_i _02080_ _00309_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13538_ _03931_ _03990_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11987__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13768__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13469_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _05592_ vssd1 vssd1
+ vccd1 vccd1 _03930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16257_ clknet_leaf_97_wb_clk_i net1739 _00245_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15208_ net1289 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16188_ clknet_leaf_115_wb_clk_i _01948_ _00176_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15139_ net1186 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18044__1544 vssd1 vssd1 vccd1 vccd1 _18044__1544/HI net1544 sky130_fd_sc_hd__conb_1
XFILLER_0_103_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09700_ net1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[21\] net945
+ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12611__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08543__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11142__A3 _07014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09631_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[23\] net953
+ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_88_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09562_ _05898_ _05900_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14092__A2 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08513_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[18\] net934
+ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09493_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\] net702 _05828_ _05832_
+ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_37_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13848__A_N net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17973__1473 vssd1 vssd1 vccd1 vccd1 _17973__1473/HI net1473 sky130_fd_sc_hd__conb_1
XFILLER_0_93_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08444_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[23\] net907 vssd1
+ vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__and3_1
XANTENNA__15223__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08375_ _04626_ _04711_ _04712_ _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__or4_2
XFILLER_0_129_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout423_A _07966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1165_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09271__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11897__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13355__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09023__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout792_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09891__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1407 net1413 vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__buf_4
Xfanout420 net422 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__clkbuf_8
Xfanout431 net434 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout442 _07962_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout453 net454 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__buf_6
XANTENNA__12521__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout464 net466 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout475 net478 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout486 _07948_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08938__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09829_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[13\] net817 net812 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__a22o_1
Xfanout497 net498 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_31_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12840_ net2298 net212 net380 vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__mux2_1
XANTENNA__14083__A2 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12094__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12771_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] net1055 net364 _03608_
+ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08837__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14510_ net1333 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__inv_2
XANTENNA__15133__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11722_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] _07798_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07915_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15490_ net1262 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09131__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08673__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ net721 _07621_ net616 _07859_ vssd1 vssd1 vccd1 vccd1 _07860_ sky130_fd_sc_hd__o211a_1
X_14441_ net1376 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__inv_2
XANTENNA__09247__C1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10277__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09798__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10604_ _06941_ _06943_ net542 vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__mux2_1
XANTENNA__13594__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17160_ clknet_leaf_22_wb_clk_i _02847_ _01143_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14372_ net1343 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11584_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] _07800_ vssd1 vssd1 vccd1
+ vccd1 _07801_ sky130_fd_sc_hd__and2_1
XANTENNA__08970__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09262__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13323_ _04477_ _03801_ _04518_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__a21o_1
X_16111_ clknet_leaf_99_wb_clk_i _01886_ _00099_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10535_ _06871_ _06872_ _06873_ _06874_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__or4_1
XFILLER_0_134_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17091_ clknet_leaf_22_wb_clk_i _02778_ _01074_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16817__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13346__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16042_ clknet_leaf_66_wb_clk_i _01836_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13254_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] _03744_ vssd1 vssd1 vccd1 vccd1
+ _03746_ sky130_fd_sc_hd__or2_1
X_10466_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[26\] net777 net748 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12205_ net1822 net269 net443 vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__mux2_1
XANTENNA__13100__B net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ net25 net837 net630 net2078 vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__a22o_1
X_10397_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\] net767 _06730_ _06736_
+ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__o22a_2
XFILLER_0_62_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10443__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09970__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12136_ net3232 net271 net454 vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__mux2_1
XANTENNA__16967__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17993_ net1493 vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__buf_2
XANTENNA__09009__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13649__A2 _07507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12067_ net2279 net205 net459 vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__mux2_1
XANTENNA__12431__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16944_ clknet_leaf_127_wb_clk_i _02631_ _00927_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_97_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08848__C _05154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09722__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11018_ _04883_ _06671_ vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_105_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16875_ clknet_leaf_0_wb_clk_i _02562_ _00858_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_26_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_105_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15826_ net1372 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14074__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13770__B _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12085__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13282__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15757_ net1401 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__inv_2
X_12969_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[117\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[125\]
+ net857 vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14708_ net1305 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15688_ net1289 vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08583__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15978__A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17427_ clknet_leaf_137_wb_clk_i _03114_ _01410_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14639_ net1225 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10187__A _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09789__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08160_ net1876 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[113\] net1052 vssd1 vssd1
+ vccd1 vccd1 _03527_ sky130_fd_sc_hd__mux2_1
XANTENNA__09976__A _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17358_ clknet_leaf_5_wb_clk_i _03045_ _01341_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16309_ clknet_leaf_75_wb_clk_i _02063_ _00292_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08091_ _04525_ _04561_ _04562_ net570 net1645 vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__a32o_1
XANTENNA__16497__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12606__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17289_ clknet_leaf_23_wb_clk_i _02976_ _01272_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10634__B _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10020__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09961__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[8\] net913 vssd1
+ vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11168__D _07507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15218__A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12341__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08758__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11465__B net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout373_A _06465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17122__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09614_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[24\] _04636_ net787
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[24\] vssd1 vssd1 vccd1 vccd1
+ _05954_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10874__A2 _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14065__A2 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09545_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[28\] net783 net754 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[28\]
+ _05871_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout540_A _05189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1282_A net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11823__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09476_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[30\] net670 net668 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[30\]
+ _05810_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_138_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08266__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08427_ net1106 net1112 net1115 net1109 vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__nor4b_4
XTAP_TAPCELL_ROW_134_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout805_A _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09886__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13576__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08358_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[30\] net821 _04647_ _04679_
+ _04683_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_24_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12516__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08289_ net1146 net1148 net1152 net1153 vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_62_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13839__C team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10825__A _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11420__S _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[18\] net962
+ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10251_ net340 vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10011__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10182_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[10\] net821 net782 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1204 net1415 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1215 net1218 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1226 net1227 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__buf_2
XANTENNA__12251__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1237 net1240 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__buf_4
X_14990_ net1284 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout250 _07842_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08507__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout1248 net1249 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__buf_4
Xfanout261 net262 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_2
Xfanout1259 net1261 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13500__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09126__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout272 net273 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_2
XANTENNA__08668__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13941_ _04218_ _04232_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__nor2_4
Xfanout283 net286 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__buf_2
Xfanout294 _07926_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_2
XANTENNA__08030__A team_01_WB.instance_to_wrap.cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_89_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16660_ clknet_leaf_128_wb_clk_i _02347_ _00643_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13872_ net160 net71 net73 vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__and3b_1
XANTENNA__08965__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15611_ net1197 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12823_ net1033 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[3\] vssd1 vssd1 vccd1
+ vccd1 _03645_ sky130_fd_sc_hd__or2_1
X_16591_ clknet_leaf_1_wb_clk_i _02278_ _00574_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_74_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15542_ net1270 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__inv_2
XANTENNA__08176__S net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12754_ net1025 _07600_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__nand2_1
XANTENNA__09483__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11705_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[10\] net717 vssd1 vssd1 vccd1
+ vccd1 _07901_ sky130_fd_sc_hd__or2_1
X_18043__1543 vssd1 vssd1 vccd1 vccd1 _18043__1543/HI net1543 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_117_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ net2299 net316 net388 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__mux2_1
X_15473_ net1293 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_144_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_144_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17212_ clknet_leaf_37_wb_clk_i _02899_ _01195_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14424_ net1361 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__inv_2
X_11636_ net616 _07846_ _07843_ _07844_ vssd1 vssd1 vccd1 vccd1 _07847_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09235__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17143_ clknet_leaf_136_wb_clk_i _02830_ _01126_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11567_ net3200 net154 team_01_WB.instance_to_wrap.cpu.K0.next_state vssd1 vssd1
+ vccd1 vccd1 _03273_ sky130_fd_sc_hd__mux2_1
X_14355_ net1364 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__inv_2
XANTENNA__12426__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10250__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11330__S _07655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13111__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10518_ net503 vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__inv_2
X_13306_ net565 _07711_ _03788_ net829 vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__a31o_1
XANTENNA__13319__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold709 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
X_17074_ clknet_leaf_134_wb_clk_i _02761_ _01057_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14286_ net1374 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11498_ net1701 net877 _07758_ _07776_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__o22a_1
XFILLER_0_81_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16025_ net1366 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13237_ net3116 net355 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1
+ vccd1 vccd1 _01913_ sky130_fd_sc_hd__a22o_1
X_10449_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[26\] net974
+ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17972__1472 vssd1 vssd1 vccd1 vccd1 _17972__1472/HI net1472 sky130_fd_sc_hd__conb_1
X_13168_ net2044 net849 net841 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[8\] vssd1
+ vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17145__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ net2709 net309 net456 vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12161__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17976_ net1476 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
X_13099_ _03719_ _03720_ _03721_ _03722_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__or4_1
Xhold1409 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16927_ clknet_leaf_25_wb_clk_i _02614_ _00910_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11285__B _07566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13781__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16858_ clknet_leaf_45_wb_clk_i _02545_ _00841_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14047__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17295__CLK clknet_leaf_143_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15809_ net1310 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__inv_2
X_16789_ clknet_leaf_122_wb_clk_i _02476_ _00772_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[24\] net676 net668 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_111_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09261_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[20\] net693 net676 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09202__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08212_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[69\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[61\]
+ net1039 vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13558__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10348__C net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09192_ net1075 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[17\] net919
+ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09226__A2 _05564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08143_ _04479_ team_01_WB.instance_to_wrap.cpu.f0.num\[15\] _04498_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\]
+ _04589_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__o221a_1
XFILLER_0_114_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12336__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout219_A _07835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10241__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08074_ _04524_ _04547_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10792__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08115__A team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1030_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1128_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09934__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13730__B2 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout490_A _07947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout588_A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12071__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 _03495_ vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[8\] net913 vssd1
+ vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold25 team_01_WB.instance_to_wrap.cpu.f0.write_data\[16\] vssd1 vssd1 vccd1 vccd1
+ net1641 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09147__D1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold36 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[30\] vssd1 vssd1 vccd1 vccd1
+ net1652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 _01828_ vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 _02077_ vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17638__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold69 net150 vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_85_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold1403_A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout922_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16662__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ _05805_ _05807_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_45_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09459_ _05784_ _05796_ _05797_ _05798_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__or4_1
XFILLER_0_93_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15411__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10258__C _06472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13549__A1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12470_ net2546 net237 net411 vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__mux2_1
XANTENNA__17018__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09217__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12754__B _07600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11421_ net327 _07733_ _07734_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12246__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10555__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10232__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14140_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[95\] _04241_ _04256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[47\]
+ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11352_ _04481_ _07680_ vssd1 vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_128_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10303_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[18\] net755 net753 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__a22o_1
X_14071_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[68\] _04247_ _04253_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__a22o_1
XANTENNA__17168__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11283_ _07188_ _07232_ _07553_ _07600_ vssd1 vssd1 vccd1 vccd1 _07623_ sky130_fd_sc_hd__or4b_1
XFILLER_0_123_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13022_ net1874 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[72\] net868 vssd1 vssd1
+ vccd1 vccd1 _02103_ sky130_fd_sc_hd__mux2_1
X_10234_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[9\] net797 net792 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__a22o_1
XANTENNA_input51_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1001 net1014 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__buf_2
Xfanout1012 net1013 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__buf_2
X_17830_ clknet_leaf_64_wb_clk_i _03506_ _01770_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[100\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_101_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11386__A team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10165_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[10\] net802 net732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[10\]
+ _06504_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_7_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10290__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1023 net1024 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16192__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1034 net1035 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__buf_2
Xfanout1045 team_01_WB.instance_to_wrap.cpu.SR1.enable vssd1 vssd1 vccd1 vccd1 net1045
+ sky130_fd_sc_hd__buf_2
Xfanout1056 team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1 vccd1
+ net1056 sky130_fd_sc_hd__buf_2
X_17761_ clknet_leaf_79_wb_clk_i _03437_ _01701_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1067 team_01_WB.instance_to_wrap.cpu.IM0.pc_enable vssd1 vssd1 vccd1 vccd1
+ net1067 sky130_fd_sc_hd__buf_2
X_14973_ net1263 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__inv_2
X_10096_ _06426_ _06430_ _06435_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__or3_4
Xfanout1078 net1096 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1089 net1096 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__clkbuf_4
X_16712_ clknet_leaf_30_wb_clk_i _02399_ _00695_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13924_ net3036 _04215_ _04216_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__o21a_1
XANTENNA__10838__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17692_ clknet_leaf_96_wb_clk_i _03376_ _01633_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14029__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_137_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12929__B net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16643_ clknet_leaf_19_wb_clk_i _02330_ _00626_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13855_ net1163 net1058 net3291 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[16\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ net2063 net641 net608 _03632_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__a22o_1
X_16574_ clknet_leaf_59_wb_clk_i _02261_ _00557_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13786_ _04158_ _04169_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10998_ net556 _05263_ _06902_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__or3_1
XANTENNA__09456__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15525_ net1210 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__inv_2
XANTENNA__09022__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12737_ net2108 net642 net606 _03585_ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a22o_1
XANTENNA__10471__B1 _06809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15456_ net1244 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12668_ net2790 net235 net387 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__mux2_1
XANTENNA__09957__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08861__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14407_ net1376 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__inv_2
XANTENNA__12156__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _07819_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\]
+ vssd1 vssd1 vccd1 vccd1 _07833_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15387_ net1180 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__inv_2
X_12599_ net2314 net245 net395 vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17126_ clknet_leaf_38_wb_clk_i _02813_ _01109_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12763__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14338_ net1371 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__inv_2
Xhold506 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10184__B net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11995__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold517 team_01_WB.instance_to_wrap.cpu.f0.write_data\[9\] vssd1 vssd1 vccd1 vccd1
+ net2133 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13776__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold528 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17057_ clknet_leaf_43_wb_clk_i _02744_ _01040_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold539 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14269_ net1321 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09916__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16008_ net1386 vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_41_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11296__A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__A1 _05570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08830_ net1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[1\] net932 vssd1
+ vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1206 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08761_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[4\] net658 _05084_ _05095_
+ _05098_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__a2111o_1
Xhold1217 team_01_WB.instance_to_wrap.cpu.f0.num\[19\] vssd1 vssd1 vccd1 vccd1 net2833
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17959_ net1459 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
Xhold1228 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2844 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1239 team_01_WB.instance_to_wrap.cpu.f0.num\[17\] vssd1 vssd1 vccd1 vccd1 net2855
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16685__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08692_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[7\] net682 _05009_ _05011_
+ _05016_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_79_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11743__B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09447__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09313_ _05649_ _05650_ _05651_ _05652_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__or4_1
XFILLER_0_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout336_A _06912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10078__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09244_ _05572_ _05581_ _05582_ _05583_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__or4_1
XANTENNA__10462__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1078_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08771__C net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09175_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[16\] net938
+ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__o21a_1
XANTENNA__12066__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13400__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17310__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout503_A _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1245_A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ _04473_ team_01_WB.instance_to_wrap.cpu.f0.num\[21\] team_01_WB.instance_to_wrap.cpu.f0.num\[17\]
+ _04477_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_47_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10765__A1 _05867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08057_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\] team_01_WB.instance_to_wrap.cpu.K0.keyvalid
+ _04523_ _04534_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1412_A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout872_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18042__1542 vssd1 vssd1 vccd1 vccd1 _18042__1542/HI net1542 sky130_fd_sc_hd__conb_1
XFILLER_0_76_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08959_ _05290_ _05291_ _05297_ _05298_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__or4_1
X_11970_ net2506 net246 net471 vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09686__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08946__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10921_ net524 _07218_ _07150_ _07040_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_58_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10852_ _06501_ _06530_ _07191_ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__or3_1
X_13640_ net983 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] _04075_ _04076_
+ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17971__1471 vssd1 vssd1 vccd1 vccd1 _17971__1471/HI net1471 sky130_fd_sc_hd__conb_1
X_10783_ _06944_ _06950_ net520 vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13571_ net980 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] _04017_ _04018_
+ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16408__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15310_ net1297 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12522_ _07793_ _07951_ net573 vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__and3_4
X_16290_ clknet_leaf_61_wb_clk_i _02044_ _00273_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[13\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_125_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08681__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15241_ net1228 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__inv_2
X_12453_ net3195 net318 net418 vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11404_ _07695_ net327 _07725_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__and3b_1
XFILLER_0_105_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12384_ net2130 net296 net426 vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__mux2_1
XANTENNA__16558__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15172_ net1239 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09610__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14123_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[14\] _04253_ _04256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[46\]
+ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__a22o_1
X_11335_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\] team_01_WB.instance_to_wrap.cpu.f0.state\[4\]
+ _04559_ _07652_ vssd1 vssd1 vccd1 vccd1 _07666_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12704__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14054_ _04236_ _04247_ _04258_ _04259_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__or4_1
X_11266_ net375 _06918_ net332 vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10732__B _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13170__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13005_ net2893 net2856 net867 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__mux2_1
X_10217_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[8\] net791 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11197_ _05529_ net332 _07536_ net370 vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__a211o_1
XANTENNA__10451__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17813_ clknet_leaf_71_wb_clk_i net2816 _01753_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[83\]
+ sky130_fd_sc_hd__dfrtp_1
X_10148_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[11\] net800 net757 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09017__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17744_ clknet_leaf_85_wb_clk_i _03420_ _01684_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14956_ net1184 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__inv_2
X_10079_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[7\] net949 vssd1
+ vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__and3_1
XANTENNA__09677__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] _04204_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__a21o_1
XANTENNA__12681__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17675_ clknet_leaf_111_wb_clk_i _03360_ _01616_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14887_ net1327 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16626_ clknet_leaf_134_wb_clk_i _02313_ _00609_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13838_ net1982 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[31\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_134_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09429__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16557_ clknet_leaf_116_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[23\]
+ _00540_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13769_ _04156_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15508_ net1313 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16488_ clknet_leaf_97_wb_clk_i _02242_ _00471_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10995__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15439_ net1218 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold303 team_01_WB.instance_to_wrap.a1.ADR_I\[26\] vssd1 vssd1 vccd1 vccd1 net1919
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold314 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
X_17109_ clknet_leaf_124_wb_clk_i _02796_ _01092_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold325 _02157_ vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12614__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18089_ net1586 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
Xhold336 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 team_01_WB.instance_to_wrap.a1.ADR_I\[19\] vssd1 vssd1 vccd1 vccd1 net1974
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[4\] net779 net746 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__a22o_1
Xhold369 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout805 _04641_ vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_6
Xfanout816 _04636_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_8
XANTENNA__09365__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09862_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[12\] net816 net770 _06196_
+ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__a211o_1
Xfanout827 net828 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout838 _03736_ vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_2
Xfanout849 net851 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_4
Xhold1003 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[63\] vssd1 vssd1 vccd1 vccd1
+ net2619 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] net730 vssd1 vssd1 vccd1 vccd1
+ _05153_ sky130_fd_sc_hd__and2_1
Xhold1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ _06129_ _06131_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__nor2_1
Xhold1025 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout286_A _07908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1036 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[47\] vssd1 vssd1 vccd1 vccd1
+ net2663 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[4\] net879 vssd1
+ vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__and3_1
Xhold1058 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1069 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[66\] vssd1 vssd1 vccd1 vccd1
+ net2685 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11473__B net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08675_ net1073 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[7\] net922 vssd1
+ vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout453_A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1195_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10683__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1362_A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout718_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08274__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09597__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09840__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09227_ _05529_ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_63_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09158_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[16\] net902
+ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08109_ _04504_ net1162 vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09089_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[13\] net914
+ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__and3_1
XANTENNA__12524__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11120_ _06313_ net334 net333 vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08303__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold870 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 _02138_ vssd1 vssd1 vccd1 vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ _07389_ _07390_ _07388_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13152__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08022__B _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ net516 _06341_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10271__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17206__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14810_ net1192 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__inv_2
X_15790_ net1316 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__inv_2
XANTENNA__09134__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1570 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[95\] vssd1 vssd1 vccd1 vccd1
+ net3186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08676__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ net1308 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__inv_2
Xhold1581 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3197 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11383__B _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11953_ net3189 net309 net476 vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__mux2_1
Xhold1592 team_01_WB.instance_to_wrap.a1.curr_state\[0\] vssd1 vssd1 vccd1 vccd1 net3208
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16230__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17460_ clknet_leaf_12_wb_clk_i _03147_ _01443_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10904_ net336 _07243_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14672_ net1377 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11884_ net2450 net281 net483 vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__mux2_1
X_16411_ clknet_leaf_67_wb_clk_i _02165_ _00394_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13623_ net982 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] _04061_ _04062_
+ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10835_ _06193_ _06218_ _07173_ _06192_ _06164_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__a311oi_4
X_17391_ clknet_leaf_142_wb_clk_i _03078_ _01374_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11218__A2 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08619__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16342_ clknet_leaf_68_wb_clk_i net2918 _00325_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08184__S net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13554_ net722 _07621_ net1066 vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__o21a_1
X_10766_ _07104_ _07105_ net522 vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__mux2_1
XANTENNA__09831__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10977__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12505_ net2169 net265 net408 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
X_16273_ clknet_leaf_68_wb_clk_i _00001_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10697_ _06941_ _06949_ net534 vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__mux2_1
X_13485_ _03850_ _03851_ _03943_ _03848_ _03847_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a311o_1
XANTENNA__09300__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18012_ net1512 vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_hd__buf_2
XANTENNA__10446__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15224_ net1176 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__inv_2
X_12436_ net2628 net241 net415 vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15155_ net1279 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12434__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ net2363 net202 net423 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__mux2_1
XANTENNA__14215__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14106_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[37\] _04230_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[117\]
+ _04392_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ _04505_ _07652_ _07654_ _07650_ vssd1 vssd1 vccd1 vccd1 _07655_ sky130_fd_sc_hd__a211o_4
X_15086_ net1282 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__inv_2
X_12298_ net2310 net210 net433 vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__mux2_1
XANTENNA__13143__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14037_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] _04265_ _04289_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ _04152_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__a221o_1
X_11249_ _07588_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09898__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11574__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15988_ net1394 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__inv_2
XANTENNA__08586__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17727_ clknet_leaf_86_wb_clk_i _03404_ _01668_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_14939_ net1195 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08460_ net1011 net885 vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__and2_2
X_17658_ clknet_leaf_90_wb_clk_i _03343_ _01599_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16609_ clknet_leaf_48_wb_clk_i _02296_ _00592_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08391_ _04724_ _04730_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12609__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17589_ clknet_leaf_80_wb_clk_i _03276_ _01548_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11513__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12957__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18041__1541 vssd1 vssd1 vccd1 vccd1 _18041__1541/HI net1541 sky130_fd_sc_hd__conb_1
XFILLER_0_50_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09210__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09012_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[9\] net939 vssd1
+ vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold100 team_01_WB.instance_to_wrap.cpu.f0.write_data\[22\] vssd1 vssd1 vccd1 vccd1
+ net1716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12344__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold111 team_01_WB.instance_to_wrap.cpu.f0.write_data\[19\] vssd1 vssd1 vccd1 vccd1
+ net1727 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold122 net85 vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold133 _03413_ vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11393__A1 _04466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17229__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold155 team_01_WB.instance_to_wrap.a1.ADR_I\[15\] vssd1 vssd1 vccd1 vccd1 net1771
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1
+ net1782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold177 _02009_ vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09338__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold188 _01973_ vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _06250_ _06253_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__nand2_1
Xhold199 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[0\] vssd1 vssd1 vccd1 vccd1 net1815
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 _04754_ vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_4
Xfanout613 net614 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_2
Xfanout624 _04628_ vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1110_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17970__1470 vssd1 vssd1 vccd1 vccd1 _17970__1470/HI net1470 sky130_fd_sc_hd__conb_1
Xfanout635 _03733_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1208_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout646 _04839_ vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__clkbuf_2
Xfanout657 _04815_ vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__buf_6
X_09845_ _06180_ _06182_ _06183_ _06184_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__or4_1
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11696__A2 _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 net669 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_8
Xfanout679 net680 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_6
XANTENNA__16253__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17379__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14095__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08269__S net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[15\] net806 net748 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13437__A3 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08727_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[5\] net693 _05054_ _05056_
+ _05062_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_94_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout835_A _03737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09889__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08658_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[10\] net698 _04978_
+ _04979_ _04990_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10120__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold246_A team_01_WB.instance_to_wrap.cpu.f0.write_data\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12519__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[15\] net692 net659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10620_ _06934_ _06959_ _06927_ _06933_ vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_137_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10551_ _06707_ net372 net544 vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09120__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10266__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13270_ net586 _03750_ _03759_ _03760_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__a31o_1
X_10482_ _06814_ _06820_ vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12221_ net2440 net314 net446 vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__mux2_1
XANTENNA__11659__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13373__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12254__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10563__A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12152_ net2297 net310 net453 vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__mux2_1
XANTENNA__09129__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11103_ net556 _06280_ net334 _07442_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16960_ clknet_leaf_32_wb_clk_i _02647_ _00943_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12083_ net2135 net279 net459 vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08968__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15911_ net1410 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__inv_2
X_11034_ net377 net341 vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__xnor2_1
X_16891_ clknet_leaf_20_wb_clk_i _02578_ _00874_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12884__A1 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13085__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15842_ net1357 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__inv_2
XANTENNA__16746__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ net1322 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__inv_2
X_12985_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[101\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[109\]
+ net857 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ clknet_leaf_23_wb_clk_i _03199_ _01495_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14724_ net1343 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11936_ net2444 net245 net475 vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__mux2_1
XANTENNA__10111__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17443_ clknet_leaf_23_wb_clk_i _03130_ _01426_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14655_ net1312 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12429__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11867_ net2621 net277 net485 vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16896__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12939__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13606_ net199 net195 _07807_ _07895_ net645 vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_67_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17374_ clknet_leaf_48_wb_clk_i _03061_ _01357_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10818_ _07156_ _07157_ net521 vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14586_ net1387 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__inv_2
XANTENNA__09265__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09804__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11798_ net2117 net211 net493 vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16325_ clknet_leaf_75_wb_clk_i net2377 _00308_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11072__B1 _07364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13537_ _03925_ _03935_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__or2_1
X_10749_ _06744_ _06747_ _06106_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16256_ clknet_leaf_96_wb_clk_i net1866 _00244_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
XANTENNA__14010__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13468_ _03926_ _03928_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15207_ net1327 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12419_ net2895 net305 net421 vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__mux2_1
X_16187_ clknet_leaf_113_wb_clk_i _01947_ _00175_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10473__A _05729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12164__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10178__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13399_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ net595 vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15138_ net1266 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__inv_2
XANTENNA__11288__B team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16276__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15069_ net1244 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12875__A1 _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09630_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[23\] net945
+ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__and3_1
XANTENNA__08543__A2 _04881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17671__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09561_ _05898_ _05900_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__nand2_1
XANTENNA__09205__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08512_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[18\] net922 vssd1
+ vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09492_ _05816_ _05819_ _05830_ _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09502__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08443_ net1010 net906 vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_1196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12339__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08374_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] net1155 vssd1 vssd1 vccd1
+ vccd1 _04714_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1060_A team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout416_A _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1158_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14001__B1 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13355__A2 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12074__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16619__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10169__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1325_A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout785_A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11118__A1 _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1408 net1413 vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__clkbuf_4
Xfanout410 _03564_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout421 net422 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_8
XANTENNA__16769__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout432 net434 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13512__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout443 _07959_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_126_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12866__A1 net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout454 _07957_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout952_A _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout465 net466 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_6
Xfanout476 net478 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08534__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09828_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[13\] net798 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__a22o_1
Xfanout487 _07947_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_6
Xfanout498 _07943_ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_6
XFILLER_0_9_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09759_ _05618_ _05731_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_100_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09495__A0 _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12770_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[19\] _07135_ net1027 vssd1 vssd1
+ vccd1 vccd1 _03608_ sky130_fd_sc_hd__mux2_1
X_11721_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[7\] net719 net615 vssd1 vssd1
+ vccd1 vccd1 _07914_ sky130_fd_sc_hd__o21a_1
XANTENNA__12249__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16149__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14440_ net1376 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__inv_2
X_11652_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[21\] net715 vssd1 vssd1 vccd1
+ vccd1 _07859_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08028__A team_01_WB.instance_to_wrap.cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10603_ net551 _06496_ _06942_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14371_ net1343 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__inv_2
XANTENNA__13594__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11583_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\]
+ _07798_ vssd1 vssd1 vccd1 vccd1 _07800_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16110_ clknet_leaf_91_wb_clk_i _01885_ _00098_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13322_ net610 _07703_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17090_ clknet_leaf_35_wb_clk_i _02777_ _01073_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10534_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[31\] net698 net679 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16041_ clknet_leaf_67_wb_clk_i _01835_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10465_ _06801_ _06802_ _06803_ _06804_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__or4_1
X_13253_ _03744_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_1310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17544__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12204_ net2931 net235 net443 vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10396_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[16\] net793 _06731_
+ _06734_ _06735_ vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__a2111o_1
X_13184_ net26 net835 net628 net1982 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12135_ net2521 net246 net451 vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17992_ net1492 vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__buf_2
XANTENNA__12712__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11109__A1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16943_ clknet_leaf_142_wb_clk_i _02630_ _00926_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12066_ net2215 net274 net461 vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18040__1540 vssd1 vssd1 vccd1 vccd1 _18040__1540/HI net1540 sky130_fd_sc_hd__conb_1
X_11017_ _07355_ _07356_ _07353_ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_105_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16874_ clknet_leaf_11_wb_clk_i _02561_ _00857_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15825_ net1321 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15756_ net1400 vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__inv_2
X_12968_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[118\] net1940 net852 vssd1 vssd1
+ vccd1 vccd1 _02157_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09486__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13282__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08864__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14707_ net1304 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__inv_2
X_11919_ net2797 net295 net481 vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15687_ net1326 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__inv_2
XANTENNA__12159__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ net357 _03673_ _03674_ net870 net2031 vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_64_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17426_ clknet_leaf_129_wb_clk_i _03113_ _01409_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14638_ net1324 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__inv_2
XANTENNA__17074__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09238__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11998__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13779__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17357_ clknet_leaf_138_wb_clk_i _03044_ _01340_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14569_ net1402 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16308_ clknet_leaf_79_wb_clk_i _02062_ _00291_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12793__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08090_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] _04524_ vssd1 vssd1 vccd1 vccd1
+ _04562_ sky130_fd_sc_hd__or2_1
X_17288_ clknet_leaf_22_wb_clk_i _02975_ _01271_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15994__A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16239_ clknet_leaf_84_wb_clk_i _01999_ _00227_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_77_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09410__B1 _04808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16911__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08104__C _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12622__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[8\] net881 vssd1
+ vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_75_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10859__A0 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout199_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10323__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09613_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[24\] net762 net752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[24\]
+ _05940_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10874__A3 _05931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout366_A _03580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09544_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[28\] net808 net752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09477__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09475_ net1071 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[30\] net893
+ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__and3_1
XANTENNA__12069__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout533_A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1275_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08426_ net1078 net926 vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_134_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13576__A2 _07231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout700_A _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08357_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[30\] net815 net794 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__a22o_1
XANTENNA__16441__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12784__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08288_ _04625_ _04626_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10825__B net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10250_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] _06589_ net624 vssd1
+ vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__mux2_1
XANTENNA__16591__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09401__B1 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10181_ _06503_ _06519_ _06520_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_37_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12532__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1205 net1211 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__buf_4
Xfanout1216 net1218 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__buf_4
XANTENNA__08949__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08311__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1227 net1236 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__clkbuf_4
Xfanout1238 net1240 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__buf_2
Xfanout240 _07870_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout251 _07904_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_2
Xfanout1249 net1269 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__clkbuf_4
Xfanout262 _07888_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_22_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08507__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13940_ _04228_ _04231_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__nand2_2
Xfanout273 _07866_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_2
XANTENNA__13500__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout284 net286 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_2
XANTENNA__11511__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08030__B _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout295 _07926_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13871_ net1617 net1168 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.next_keyvalid
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15610_ net1192 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
X_12822_ net1033 net322 vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13264__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16590_ clknet_leaf_8_wb_clk_i _02277_ _00573_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_16_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08684__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15541_ net1225 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__inv_2
XANTENNA__11275__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12753_ net2678 net639 net606 _03596_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__a22o_1
XANTENNA__14983__A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11704_ net2119 net227 net501 vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15472_ net1226 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__inv_2
X_12684_ net2404 net318 net388 vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__mux2_1
XANTENNA__08981__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17211_ clknet_leaf_19_wb_clk_i _02898_ _01194_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ net1361 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ _07818_ _07845_ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__or2_1
XANTENNA__12707__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11611__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17142_ clknet_leaf_141_wb_clk_i _02829_ _01125_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14354_ net1371 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11566_ team_01_WB.instance_to_wrap.cpu.K0.count\[0\] team_01_WB.instance_to_wrap.cpu.K0.count\[1\]
+ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__nand2b_1
XFILLER_0_25_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10250__A1 _06589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13305_ _04473_ _07709_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13111__B net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10517_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] net625 _06855_ _06856_
+ vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__a22o_2
X_17073_ clknet_leaf_14_wb_clk_i _02760_ _01056_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14285_ net1374 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11497_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[14\] _07756_ vssd1 vssd1 vccd1
+ vccd1 _07776_ sky130_fd_sc_hd__and2_1
XANTENNA__10454__C net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_113_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16024_ net1351 vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__inv_2
X_13236_ team_01_WB.instance_to_wrap.cpu.f0.num\[14\] net356 net352 net2660 vssd1
+ vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a22o_1
X_10448_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[26\] net946
+ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15319__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12442__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ net2071 net850 net842 net1955 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__a22o_1
X_10379_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[16\] net790 net750 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12118_ net1977 net294 net456 vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__mux2_1
XANTENNA__08859__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17975_ net1475 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
X_13098_ net43 net42 net45 net44 vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__or4_2
X_16926_ clknet_leaf_44_wb_clk_i _02613_ _00909_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12049_ net2311 net304 net463 vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10305__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16314__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16857_ clknet_leaf_51_wb_clk_i _02544_ _00840_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11582__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15808_ net1342 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__inv_2
X_16788_ clknet_leaf_12_wb_clk_i _02475_ _00771_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11266__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15739_ net1184 vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09260_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[20\] net689 net679 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08211_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[70\] net2512 net1042 vssd1 vssd1
+ vccd1 vccd1 _03476_ sky130_fd_sc_hd__mux2_1
X_17409_ clknet_leaf_48_wb_clk_i _03096_ _01392_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13558__A2 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09191_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[17\] net934 vssd1
+ vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__and3_1
XANTENNA__12617__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12766__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08142_ _04474_ team_01_WB.instance_to_wrap.cpu.f0.num\[20\] team_01_WB.instance_to_wrap.cpu.f0.num\[7\]
+ _04486_ _04597_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__o221a_1
XFILLER_0_132_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08073_ _04525_ _04548_ _04549_ net569 team_01_WB.instance_to_wrap.cpu.f0.write_data\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13191__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12352__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1023_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__B2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[8\] net675 _05312_ _05313_
+ _05314_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_122_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout483_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold15 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[28\] vssd1 vssd1 vccd1 vccd1
+ net1631 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold26 _03552_ vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 team_01_WB.instance_to_wrap.cpu.f0.write_data\[31\] vssd1 vssd1 vccd1 vccd1
+ net1653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[83\] vssd1 vssd1 vccd1 vccd1 net1664
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold59 team_01_WB.instance_to_wrap.cpu.f0.write_data\[30\] vssd1 vssd1 vccd1 vccd1
+ net1675 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07970__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout650_A _04823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1392_A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_A _04682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13246__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09527_ _05865_ _05866_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] net625
+ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout915_A net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09458_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[29\] _04766_ net678
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[29\] vssd1 vssd1 vccd1 vccd1
+ _05798_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09870__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16957__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13549__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08409_ _04738_ _04745_ _04736_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__and3b_1
XFILLER_0_53_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12527__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ net599 _05726_ _05728_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_136_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12757__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11420_ team_01_WB.instance_to_wrap.cpu.f0.i\[16\] _07704_ _07700_ vssd1 vssd1 vccd1
+ vccd1 _07734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09622__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08306__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10555__B net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11351_ _04482_ _07678_ vssd1 vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_39_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10274__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10302_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[18\] net772 net760 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14070_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[12\] _04226_ _04256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[44\]
+ _04357_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13866__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11282_ _07088_ _07154_ net278 _07589_ vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__or4bb_1
X_13021_ net3140 net3081 net866 vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__mux2_1
XANTENNA__08728__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[9\] net801 _04649_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__a22o_1
XANTENNA__12262__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09137__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[10\] net965
+ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_89_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1002 net1004 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_7_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input44_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11386__B net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08679__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1013 net1014 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1024 _04490_ vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_8
XANTENNA__14978__A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__clkbuf_4
Xfanout1046 net1049 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17760_ clknet_leaf_75_wb_clk_i net1780 _01700_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14972_ net1172 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__inv_2
X_10095_ _06431_ _06432_ _06433_ _06434_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__or4_1
Xfanout1057 team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1 vccd1
+ net1057 sky130_fd_sc_hd__buf_2
XANTENNA__08976__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1068 team_01_WB.instance_to_wrap.cpu.IM0.pc_enable vssd1 vssd1 vccd1 vccd1
+ net1068 sky130_fd_sc_hd__clkbuf_4
Xfanout1079 net1089 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_2
X_13923_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\] _04215_ net572 vssd1
+ vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__a21boi_1
X_16711_ clknet_leaf_122_wb_clk_i _02398_ _00694_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17691_ clknet_leaf_93_wb_clk_i _03375_ _01632_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_57_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16487__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08361__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11606__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16642_ clknet_leaf_34_wb_clk_i _02329_ _00625_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17732__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13854_ net1164 net1059 net3287 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[15\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13237__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12805_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] net1056 net365 _03631_
+ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__a22o_1
X_16573_ clknet_leaf_58_wb_clk_i _02260_ _00556_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_18_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13785_ _04156_ _01836_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__nand2_1
XANTENNA__09303__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10997_ _06915_ _07325_ _07336_ net552 _07335_ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__o221a_1
XANTENNA__13642__D1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15524_ net1191 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__inv_2
XANTENNA__10449__C net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12736_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] net1054 net363 _03584_
+ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09861__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17882__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10471__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15455_ net1256 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12667_ net2088 net240 net387 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__mux2_1
XANTENNA__12437__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14406_ net1339 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__inv_2
X_11618_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[28\] _07088_ net716 vssd1 vssd1
+ vccd1 vccd1 _07832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15386_ net1190 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__inv_2
XANTENNA__09613__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12598_ net2940 net201 net395 vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17125_ clknet_leaf_31_wb_clk_i _02812_ _01108_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08967__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14337_ net1370 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17112__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11549_ net1969 net1160 vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold507 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold518 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11971__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17056_ clknet_leaf_33_wb_clk_i _02743_ _01039_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold529 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14268_ net1317 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__inv_2
XANTENNA__13173__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16007_ net1386 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ net3147 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[31\] vssd1 vssd1
+ vccd1 vccd1 _01931_ sky130_fd_sc_hd__a22o_1
XANTENNA__11577__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13712__A2 _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12172__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14199_ _04156_ _01836_ _04181_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10526__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12920__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11296__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17262__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1207 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08760_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[4\] net648 _05077_ _05080_
+ _05091_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__a2111o_1
Xhold1218 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2834 sky130_fd_sc_hd__dlygate4sd3_1
X_17958_ net1458 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
XANTENNA__08886__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_81_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1229 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2845 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09144__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16909_ clknet_leaf_140_wb_clk_i _02596_ _00892_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_08691_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[7\] net671 _05012_ _05018_
+ _05020_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__a2111o_1
X_17889_ net107 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_10_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11516__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08352__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09213__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09312_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[22\] net685 _05632_
+ _05634_ _05635_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_48_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09510__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[21\] net679 net663 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12347__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout231_A net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09174_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[16\] net658 _05511_
+ _05512_ _05513_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18114__1593 vssd1 vssd1 vccd1 vccd1 _18114__1593/HI net1593 sky130_fd_sc_hd__conb_1
XANTENNA__13400__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08958__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ _04472_ team_01_WB.instance_to_wrap.cpu.f0.num\[23\] team_01_WB.instance_to_wrap.cpu.f0.num\[19\]
+ _04475_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__o22ai_1
XANTENNA_fanout1140_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1238_A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11962__A1 _07831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10765__A2 _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08056_ _04530_ _04531_ _04533_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__or3_2
XANTENNA__09883__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout698_A _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13164__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12082__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1405_A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout865_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[6\] net667 _05268_ _05270_
+ _05287_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__a2111o_1
X_08889_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[2\] net932 vssd1
+ vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10920_ net371 _07257_ _07259_ net337 net324 vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10851_ _06601_ _07189_ _06532_ _06594_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__a211oi_2
XANTENNA__09123__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10269__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13570_ net722 _07251_ net1066 vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__o21a_1
XANTENNA__09843__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10782_ net553 _07121_ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12521_ net2707 net291 net408 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
XANTENNA__12257__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17135__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15240_ net1275 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12452_ net2145 net308 net418 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11403_ _04471_ _07713_ vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15171_ net1188 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__inv_2
X_12383_ net2113 net299 net426 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14122_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[14\] _04226_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[110\]
+ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__a221o_1
X_11334_ _07665_ net1683 _07655_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17285__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13155__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14053_ _04224_ _04238_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11265_ _06922_ _06930_ _07071_ _07603_ _07604_ vssd1 vssd1 vccd1 vccd1 _07605_ sky130_fd_sc_hd__a32o_1
XANTENNA__10508__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ net2986 net2817 net857 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__mux2_1
X_10216_ _06534_ _06553_ _06554_ _06555_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__or4_1
XANTENNA__09374__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11196_ net335 net337 _07362_ vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17812_ clknet_leaf_66_wb_clk_i net2569 _01752_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[82\]
+ sky130_fd_sc_hd__dfrtp_1
X_10147_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[11\] net817 net739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[11\]
+ _06474_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__a221o_1
XANTENNA__13458__A1 _03914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17743_ clknet_leaf_65_wb_clk_i _03419_ _01683_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_14955_ net1295 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10078_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[7\] net954 vssd1
+ vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11336__S _07655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13906_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] _04204_ _04205_ vssd1
+ vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__o21a_1
X_14886_ net1299 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__inv_2
XANTENNA__10141__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17674_ clknet_leaf_111_wb_clk_i _03359_ _01615_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16625_ clknet_leaf_17_wb_clk_i _02312_ _00608_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10692__A1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13837_ net2078 net834 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[30\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_76_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13615__D1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16556_ clknet_leaf_117_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[22\]
+ _00539_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13768_ net1170 _04155_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__nand2_1
XANTENNA__09834__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15507_ net1281 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__inv_2
X_12719_ net3071 net291 net384 vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__mux2_1
X_16487_ clknet_leaf_96_wb_clk_i _02241_ _00470_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12167__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13699_ net1881 _04106_ _04120_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[10\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15438_ net1283 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15369_ net1231 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10747__A2 _07065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold304 _02024_ vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17108_ clknet_leaf_13_wb_clk_i _02795_ _01091_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold315 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18088_ net637 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold326 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13146__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09930_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[4\] net740 net769 vssd1
+ vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__a21o_1
X_17039_ clknet_leaf_143_wb_clk_i _02726_ _01022_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold359 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[21\] vssd1 vssd1 vccd1 vccd1
+ net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11100__A _06921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout806 _04641_ vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__buf_4
Xfanout817 net818 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_8
X_09861_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[12\] net820 net783 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__a22o_1
Xfanout828 _04579_ vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09208__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11172__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout839 net840 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_4
X_08812_ net602 _05150_ _05116_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a21o_1
XANTENNA__12630__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09792_ _06129_ _06131_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__nand2_1
Xhold1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13449__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10380__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1026 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1037 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[4\] net913 vssd1
+ vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__and3_1
XANTENNA__09505__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1048 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08674_ net1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[7\] net896 vssd1
+ vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10683__A1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16032__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1090_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17158__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13606__D1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_A _07959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1188_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15242__A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13621__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08782__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12077__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout613_A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1355_A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09226_ net598 _05564_ _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_31_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09157_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[16\] net888
+ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08108_ _04504_ net1162 vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09088_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[13\] net925
+ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout982_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13137__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08039_ net1641 net568 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1
+ vccd1 vccd1 _03552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold860 team_01_WB.instance_to_wrap.a1.ADR_I\[3\] vssd1 vssd1 vccd1 vccd1 net2476
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08303__B net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold871 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[71\] vssd1 vssd1 vccd1 vccd1
+ net2498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11050_ net520 _06339_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__nand2_1
Xhold893 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09356__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__C _04810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10001_ net550 net542 net561 vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12540__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09108__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14101__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14040__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1560 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[33\] vssd1 vssd1 vccd1 vccd1
+ net3176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1571 _03501_ vssd1 vssd1 vccd1 vccd1 net3187 sky130_fd_sc_hd__dlygate4sd3_1
X_14740_ net1308 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__inv_2
X_11952_ net2268 net294 net476 vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1582 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1593 team_01_WB.instance_to_wrap.a1.ADR_I\[10\] vssd1 vssd1 vccd1 vccd1 net3209
+ sky130_fd_sc_hd__dlygate4sd3_1
X_10903_ _04883_ _06672_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__nor2_1
X_14671_ net1355 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__inv_2
X_11883_ net2748 net304 net484 vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16410_ clknet_leaf_62_wb_clk_i _02164_ _00393_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13622_ net723 _07531_ net1068 vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_120_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10834_ _06194_ _07173_ _06599_ _06164_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__o211a_1
X_17390_ clknet_leaf_10_wb_clk_i _03077_ _01373_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16341_ clknet_leaf_74_wb_clk_i _02095_ _00324_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_13553_ net185 _04002_ _04003_ net725 vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__a211o_1
X_10765_ _04706_ _05867_ _05898_ _06779_ net549 net540 vssd1 vssd1 vccd1 vccd1 _07105_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__10977__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12504_ net2064 net268 net407 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
X_16272_ clknet_leaf_68_wb_clk_i _00000_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13484_ _03848_ _03944_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__or2_1
X_10696_ _06936_ _06943_ net533 vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18011_ net1511 vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_hd__buf_2
XFILLER_0_129_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15223_ net1199 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12435_ net2971 net271 net416 vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__mux2_1
XANTENNA__12715__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15154_ net1232 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09595__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12366_ net1948 net206 net423 vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14105_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[37\] _04221_ _04260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[61\]
+ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13128__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11317_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] _04506_ team_01_WB.instance_to_wrap.cpu.f0.state\[8\]
+ _04524_ _00019_ vssd1 vssd1 vccd1 vccd1 _07654_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15085_ net1210 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12297_ net2012 net249 net433 vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__mux2_1
XANTENNA_output75_A net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14036_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[58\] _04260_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[18\]
+ _04313_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__a221o_1
XANTENNA__09347__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11248_ _07555_ _07580_ _07586_ _07587_ vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_43_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08555__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12450__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ _06903_ _07065_ _07518_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__a21o_1
XANTENNA__10362__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08867__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11574__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15987_ net1399 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17726_ clknet_leaf_87_wb_clk_i _03403_ _01667_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_19_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17300__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10114__B1 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14938_ net1187 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17657_ clknet_leaf_120_wb_clk_i _03342_ _01598_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14869_ net1221 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
XANTENNA__11590__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15062__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16608_ clknet_leaf_33_wb_clk_i _02295_ _00591_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_08390_ _04708_ _04717_ _04726_ net712 vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__nor4_1
XANTENNA__09807__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17588_ clknet_leaf_80_wb_clk_i _03275_ _01547_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09698__C net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13603__A1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09060__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17450__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16539_ clknet_leaf_90_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[5\]
+ _00522_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11090__A1 _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09011_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[9\] net932 vssd1
+ vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12625__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13310__A team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold101 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[6\] vssd1 vssd1 vccd1 vccd1 net1717
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09586__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold112 team_01_WB.instance_to_wrap.a1.ADR_I\[7\] vssd1 vssd1 vccd1 vccd1 net1728
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold123 _02017_ vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13119__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 team_01_WB.instance_to_wrap.cpu.f0.read_i vssd1 vssd1 vccd1 vccd1 net1750
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold145 net151 vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold156 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] vssd1 vssd1 vccd1 vccd1
+ net1772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[16\] vssd1 vssd1 vccd1 vccd1
+ net1783 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _05076_ _06252_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__xor2_1
XANTENNA__09338__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold178 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[11\] vssd1 vssd1 vccd1 vccd1
+ net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[95\] vssd1 vssd1 vccd1 vccd1
+ net1805 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _04754_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout614 _07636_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout396_A _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout625 net626 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 net638 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09844_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[13\] net788 net760 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__a22o_1
Xfanout647 _04825_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12360__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout658 _04815_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1103_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout669 _04801_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__buf_6
XANTENNA__08777__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09775_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[15\] net789 net776 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[5\] net661 _05044_ _05047_
+ _05052_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10105__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08849__A1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16548__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[10\] net667 _04972_
+ _04974_ _04985_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_1_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11704__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08588_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[15\] net668 net656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10408__A1 _06598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16698__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15700__A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11005__A _05729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ _06888_ _06889_ net538 vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09209_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[17\] net924
+ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12535__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10481_ _06781_ _06815_ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12220_ net2460 net318 net446 vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09577__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08314__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10563__B _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12151_ net1823 net295 net452 vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11102_ net557 net333 _07396_ net338 net371 vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_4_5__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09329__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12082_ net2885 net303 net460 vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__mux2_1
Xhold690 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15910_ net1393 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__inv_2
X_11033_ _07368_ _07371_ _07372_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12270__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17323__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16890_ clknet_leaf_46_wb_clk_i _02577_ _00873_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08687__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15841_ net1357 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_138_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_138_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_107_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ net2688 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[110\] net852 vssd1 vssd1
+ vccd1 vccd1 _02141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15772_ net1320 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1390 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[4\] vssd1 vssd1 vccd1 vccd1
+ net3006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17511_ clknet_leaf_16_wb_clk_i _03198_ _01494_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14723_ net1349 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__inv_2
X_11935_ net2266 net202 net475 vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17442_ clknet_leaf_35_wb_clk_i _03129_ _01425_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14654_ net1250 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__inv_2
X_11866_ net2347 net211 net485 vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13605_ _04029_ _04046_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__nor2_1
X_10817_ net512 net511 _06779_ _06811_ net549 net536 vssd1 vssd1 vccd1 vccd1 _07157_
+ sky130_fd_sc_hd__mux4_1
X_17373_ clknet_leaf_40_wb_clk_i _03060_ _01356_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14585_ net1402 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__inv_2
X_11797_ net2618 net249 net492 vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16324_ clknet_leaf_76_wb_clk_i net2346 _00307_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13536_ net980 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _03988_ _03989_
+ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10748_ net562 _06825_ _07057_ _07087_ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__a31o_2
XFILLER_0_83_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16255_ clknet_leaf_95_wb_clk_i net1763 _00243_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12445__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13467_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] _05655_ vssd1 vssd1
+ vccd1 vccd1 _03928_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10679_ net563 _06829_ _06962_ _07018_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__a31o_2
XANTENNA__10754__A _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15206_ net1290 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12418_ net2903 net309 net420 vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16186_ clknet_leaf_107_wb_clk_i _01946_ _00174_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13398_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] _05495_ vssd1 vssd1
+ vccd1 vccd1 _03859_ sky130_fd_sc_hd__and2_1
X_15137_ net1248 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12349_ net2434 net282 net427 vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15068_ net1173 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14019_ net1670 net605 _04309_ net1169 vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11585__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12180__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_65_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10886__A1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09560_ _05760_ _05781_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_88_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08511_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[18\] net910
+ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__and3_1
X_17709_ clknet_leaf_103_wb_clk_i _03393_ _01650_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09491_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[30\] net696 net675 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[30\]
+ _05821_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16840__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08442_ net1106 net1109 net1112 net1114 vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__and4_2
XFILLER_0_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08373_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__or2_2
XFILLER_0_92_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12355__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1053_A team_01_WB.instance_to_wrap.cpu.SR1.enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16220__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1220_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07973__A team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09891__C _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout680_A _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout400 _03566_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1409 net1413 vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__buf_4
XANTENNA__12315__A1 _07912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout411 _03563_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_8
Xfanout422 _03561_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12090__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout433 net434 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_54_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout444 _07959_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_4
Xfanout455 _07956_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_8
XANTENNA__16370__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout466 _07954_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_8
X_09827_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[13\] net779 net778 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[13\]
+ _06166_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout477 net478 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout488 _07947_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout499 _07795_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout945_A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09758_ _06096_ _06097_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] net625
+ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_9_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08709_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[5\] net908 vssd1
+ vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__and3_1
X_09689_ _06025_ _06026_ _06027_ _06028_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__or4_1
XANTENNA__13291__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11720_ net718 _07308_ vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10558__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11651_ net2096 net203 net499 vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__mux2_1
XANTENNA__09131__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10277__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08028__B _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10602_ net551 _06526_ vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__nor2_1
XANTENNA__15430__A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09798__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14370_ net1344 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__inv_2
XANTENNA__13869__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11582_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] _07798_ vssd1 vssd1 vccd1
+ vccd1 _07799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08970__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13321_ net1854 net828 _03799_ _03800_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10801__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10533_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[31\] net657 net706 vssd1
+ vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12265__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16040_ clknet_leaf_68_wb_clk_i _01834_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13252_ net610 _07710_ net1063 vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_111_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input74_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[26\] net758 _06789_ _06790_
+ _06792_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11389__B _07696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12203_ net2872 net239 net443 vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13183_ net1164 net838 team_01_WB.instance_to_wrap.a1.prev_BUSY_O vssd1 vssd1 vccd1
+ vccd1 _03739_ sky130_fd_sc_hd__or3b_1
X_10395_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[16\] net819 net778 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12134_ net3159 net202 net451 vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__mux2_1
XANTENNA__09970__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17991_ net1491 vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_27_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16713__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16942_ clknet_leaf_8_wb_clk_i _02629_ _00925_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12065_ net3141 net209 net461 vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_109_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11016_ _05618_ net507 vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__xor2_1
XANTENNA__09722__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16873_ clknet_leaf_9_wb_clk_i _02560_ _00856_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15824_ net1322 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__inv_2
XANTENNA__16863__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09603__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12967_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[119\] net1967 net862 vssd1 vssd1
+ vccd1 vccd1 _02158_ sky130_fd_sc_hd__mux2_1
X_15755_ net1400 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ net2902 net298 net482 vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__mux2_1
X_14706_ net1316 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__inv_2
X_15686_ net1326 vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__inv_2
XANTENNA__17219__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12898_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[23\] net1030 vssd1 vssd1 vccd1
+ vccd1 _03674_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_64_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17425_ clknet_leaf_15_wb_clk_i _03112_ _01408_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11849_ net2912 net285 net490 vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__mux2_1
X_14637_ net1270 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11045__A1 _05189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14568_ net1384 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__inv_2
X_17356_ clknet_leaf_131_wb_clk_i _03043_ _01339_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_35_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12793__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16307_ clknet_leaf_65_wb_clk_i net1626 _00290_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12175__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13990__B1 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13519_ net980 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _03974_ _03975_
+ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14499_ net1407 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17369__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17287_ clknet_leaf_15_wb_clk_i _02974_ _01270_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16238_ clknet_leaf_84_wb_clk_i _01998_ _00226_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_77_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16169_ clknet_leaf_100_wb_clk_i _00011_ _00157_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_58_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16393__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10020__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08991_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[8\] net672 _05328_ _05329_
+ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__09961__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10859__A1 _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09612_ _05949_ _05950_ _05951_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_30_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09543_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[28\] net748 _05872_ _05874_
+ _05881_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_92_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11462__B1_N net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout359_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10087__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09474_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[30\] net889
+ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08425_ net1109 net1113 net1114 net1106 vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_47_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1170_A _00026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout526_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15250__A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1268_A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08356_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[30\] net782 net756 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09886__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08790__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12784__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12085__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08287_ _04625_ _04626_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16736__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout895_A _04793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11002__B net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10547__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10011__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10180_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[10\] net788 net755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1206 net1211 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1217 net1218 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__buf_2
XANTENNA__16886__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1228 net1231 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__buf_4
Xfanout230 _07900_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08311__B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout241 _07870_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
XANTENNA__09165__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1239 net1240 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__buf_4
Xfanout252 _07904_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_1
XANTENNA__11282__C_N net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout263 net266 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
XANTENNA__09126__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout274 net277 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_2
Xfanout285 net286 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_2
Xfanout296 _07926_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_2
X_13870_ net1164 net1059 net3282 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[31\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__16116__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08965__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ net2180 net640 net607 _03643_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12752_ net364 _03594_ _03595_ net1055 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__a32o_1
XFILLER_0_69_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15540_ net1324 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11703_ net612 _07806_ _07899_ _07898_ vssd1 vssd1 vccd1 vccd1 _07900_ sky130_fd_sc_hd__a31o_4
X_15471_ net1217 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12683_ net2046 net307 net388 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__mux2_1
XANTENNA__16266__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08691__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ clknet_leaf_59_wb_clk_i _02897_ _01193_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ net1348 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__inv_2
XANTENNA__17511__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11634_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _07817_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\]
+ vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14353_ net1371 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__inv_2
XANTENNA__12775__B2 _03611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17141_ clknet_leaf_122_wb_clk_i _02828_ _01124_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11565_ net3210 net155 team_01_WB.instance_to_wrap.cpu.K0.next_state vssd1 vssd1
+ vccd1 vccd1 _03274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10921__A1_N net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10786__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13304_ _07686_ _07711_ _03786_ net586 vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__o211a_1
X_10516_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\] net764 net621 vssd1
+ vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17072_ clknet_leaf_15_wb_clk_i _02759_ _01055_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14284_ net1374 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__inv_2
X_11496_ net368 _07775_ net1676 net876 vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_134_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16023_ net1357 vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__inv_2
X_13235_ net3230 net355 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1
+ vccd1 vccd1 _01915_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10447_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[26\] net950
+ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__and3_1
XANTENNA__10538__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13166_ net1852 net849 net841 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[10\] vssd1
+ vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10378_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[16\] net812 net742 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[16\]
+ _06716_ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__a221o_1
X_12117_ net2110 net298 net458 vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__mux2_1
X_17974_ net1474 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
X_13097_ net70 net69 net41 net40 vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__or4_1
XFILLER_0_100_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12048_ net2934 net283 net465 vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__mux2_1
X_16925_ clknet_leaf_49_wb_clk_i _02612_ _00908_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11502__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16856_ clknet_leaf_29_wb_clk_i _02543_ _00839_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17041__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15807_ net1352 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16787_ clknet_leaf_129_wb_clk_i _02474_ _00770_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13999_ _04238_ _04242_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__nor2_1
XANTENNA__16609__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11266__A1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15738_ net1190 vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15669_ net1221 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__inv_2
XANTENNA__17191__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[71\] net3250 net1048 vssd1 vssd1
+ vccd1 vccd1 _03477_ sky130_fd_sc_hd__mux2_1
XANTENNA__11802__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17408_ clknet_leaf_30_wb_clk_i _03095_ _01391_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09190_ net1150 net619 net593 vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16759__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12766__B2 _03605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08141_ _04472_ team_01_WB.instance_to_wrap.cpu.f0.num\[23\] team_01_WB.instance_to_wrap.cpu.f0.num\[20\]
+ _04474_ _04593_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__a221o_1
X_17339_ clknet_leaf_50_wb_clk_i _03026_ _01322_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10777__A0 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10241__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08072_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] _04524_ vssd1 vssd1 vccd1 vccd1
+ _04549_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12633__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10529__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09395__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09934__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09508__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11757__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10544__A3 _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08974_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[8\] net909 vssd1
+ vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1016_A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16139__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold16 team_01_WB.instance_to_wrap.cpu.DM0.state\[1\] vssd1 vssd1 vccd1 vccd1 net1632
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold27 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[123\] vssd1 vssd1 vccd1 vccd1
+ net1643 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14140__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold38 _01832_ vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 _02122_ vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08785__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16289__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout643_A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1385_A net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\] net765 net621 vssd1
+ vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09457_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[29\] net693 net661 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout908_A _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ _04738_ _04746_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__or2_2
XFILLER_0_136_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09388_ net601 _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_95_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17684__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12757__B2 _03599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08339_ net1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[30\] net959
+ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09622__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08306__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10232__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11350_ _04482_ _07678_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _06639_ _06640_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12543__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11281_ net562 _07612_ _07613_ _07620_ vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__a31o_2
XFILLER_0_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13020_ net2685 net2608 net859 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__mux2_1
XANTENNA__09386__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[9\] net809 net737 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[9\]
+ _06570_ vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__a221o_1
XANTENNA__09925__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_5_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11732__A2 _07507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10163_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[10\] net791 net778 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__a22o_1
Xfanout1003 net1004 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_89_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1014 _04490_ vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10290__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17064__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1025 net1026 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_4
Xfanout1036 team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1 vccd1
+ net1036 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input37_A gpio_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 net1049 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__clkbuf_4
X_14971_ net1179 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__inv_2
X_10094_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[7\] net800 net750 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__a22o_1
Xfanout1058 net1059 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__clkbuf_2
Xfanout1069 net1070 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__clkbuf_2
X_16710_ clknet_leaf_38_wb_clk_i _02397_ _00693_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13922_ _04215_ net572 _04214_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__and3b_1
XANTENNA__11496__B2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17690_ clknet_leaf_94_wb_clk_i _03374_ _01631_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_57_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09153__A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16641_ clknet_leaf_42_wb_clk_i _02328_ _00624_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13853_ net1166 net1060 net2343 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[14\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__10299__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12804_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[8\] _07290_ net1033 vssd1 vssd1
+ vccd1 vccd1 _03631_ sky130_fd_sc_hd__mux2_1
X_16572_ clknet_leaf_59_wb_clk_i _02259_ _00555_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_13784_ _04162_ _04164_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08992__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10996_ _06398_ net334 net333 vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16901__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15523_ net1176 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12735_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[30\] _07019_ net1025 vssd1 vssd1
+ vccd1 vccd1 _03584_ sky130_fd_sc_hd__mux2_1
XANTENNA__12718__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11622__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12666_ net2929 net271 net389 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15454_ net1252 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12748__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14405_ net1333 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__inv_2
X_11617_ net2200 net220 net500 vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12597_ net2783 net207 net395 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__mux2_1
X_15385_ net1258 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17124_ clknet_leaf_55_wb_clk_i _02811_ _01107_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11548_ net1935 net1160 vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__and2_1
X_14336_ net1370 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold508 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12453__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14267_ net1323 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17055_ clknet_leaf_7_wb_clk_i _02742_ _01038_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold519 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
X_11479_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[23\] net579 vssd1 vssd1 vccd1
+ vccd1 _07767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09377__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13218_ team_01_WB.instance_to_wrap.cpu.f0.state\[6\] _03740_ vssd1 vssd1 vccd1 vccd1
+ _03742_ sky130_fd_sc_hd__nor2_1
X_16006_ net1358 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__inv_2
XANTENNA__09916__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11577__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14198_ net1734 _04462_ _04463_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12920__A1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13149_ net127 net845 net839 net1859 vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14122__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17957_ net1457 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
Xhold1208 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1219 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2835 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16431__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11593__A _07809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16908_ clknet_leaf_133_wb_clk_i _02595_ _00891_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_08690_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[7\] net662 _05008_ _05013_
+ _05026_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__a2111o_1
X_17888_ net107 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16839_ clknet_leaf_123_wb_clk_i _02526_ _00822_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10002__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13633__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09311_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[22\] net666 _05622_
+ _05625_ _05638_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_53_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12628__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08655__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09242_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[21\] net900
+ net657 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[21\] vssd1 vssd1 vccd1
+ vccd1 _05582_ sky130_fd_sc_hd__a32o_1
XANTENNA__10462__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12739__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09173_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[16\] net920
+ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08124_ _04481_ team_01_WB.instance_to_wrap.cpu.f0.num\[13\] team_01_WB.instance_to_wrap.cpu.f0.num\[12\]
+ _04482_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__o22a_1
XANTENNA__10214__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11411__A1 _07701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10765__A3 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08055_ _04527_ _04532_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__nor2_1
XANTENNA__12363__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1133_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09368__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12911__A1 _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1300_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14113__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__A team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08957_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[6\] net699 _05271_ _05282_
+ net708 vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout760_A _04674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08888_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[2\] net898 vssd1
+ vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11008__A _05707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ _06601_ _07189_ _06594_ vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09509_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[29\] net950
+ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__and3_1
XANTENNA__12538__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10781_ net529 _06967_ _07120_ _07119_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12520_ net2500 net314 net410 vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XANTENNA__08317__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12451_ net3033 net310 net417 vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11402_ net327 _07723_ _07724_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__and3_1
X_15170_ net1268 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__inv_2
X_12382_ net1897 net281 net425 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14121_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[94\] _04240_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[78\]
+ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11333_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] net1162 _04555_ _07652_ vssd1
+ vssd1 vccd1 vccd1 _07665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12273__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14054__A _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10582__A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09359__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14052_ _04334_ _04336_ _04338_ _04340_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__or4_1
XFILLER_0_127_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11264_ net524 _07300_ net556 vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__a21oi_1
X_13003_ net1664 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[91\] net864 vssd1 vssd1
+ vccd1 vccd1 _02122_ sky130_fd_sc_hd__mux2_1
X_10215_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[8\] net732 _06538_ _06542_
+ _06545_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08031__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11195_ net329 _07534_ vssd1 vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__and2_1
X_17811_ clknet_leaf_70_wb_clk_i _03487_ _01751_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14104__B1 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10146_ _06475_ _06478_ _06480_ _06485_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__or4_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11617__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17742_ clknet_leaf_86_wb_clk_i _03418_ _01682_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_14954_ net1279 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__inv_2
X_10077_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[7\] net967 vssd1
+ vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__and3_1
X_13905_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] _04204_ net571 vssd1
+ vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_76_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17673_ clknet_leaf_119_wb_clk_i _03358_ _01614_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14885_ net1205 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16624_ clknet_leaf_124_wb_clk_i _02311_ _00607_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13836_ net1851 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[29\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16555_ clknet_leaf_116_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[21\]
+ _00538_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13767_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[4\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ net604 vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__mux2_1
X_10979_ _06438_ net373 net340 _06562_ net552 net534 vssd1 vssd1 vccd1 vccd1 _07319_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12448__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15506_ net1235 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12718_ net2675 net315 net386 vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__mux2_1
XANTENNA__11641__B2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16486_ clknet_leaf_95_wb_clk_i _02240_ _00469_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13698_ team_01_WB.instance_to_wrap.cpu.c0.count\[10\] _04106_ _04119_ vssd1 vssd1
+ vccd1 vccd1 _04120_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15437_ net1215 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__inv_2
X_12649_ net2323 net313 net392 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10195__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15368_ net1275 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_68_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17107_ clknet_leaf_137_wb_clk_i _02794_ _01090_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11588__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12183__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold305 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1
+ net1921 sky130_fd_sc_hd__dlygate4sd3_1
X_14319_ net1178 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__inv_2
XANTENNA__10492__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold316 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
X_18087_ net637 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15299_ net1188 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold327 net121 vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold338 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold349 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
X_17038_ clknet_leaf_8_wb_clk_i _02725_ _01021_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout807 net810 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__buf_6
X_09860_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[12\] net773 _06195_
+ _06199_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__a211o_1
Xfanout818 _04634_ vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__buf_8
Xfanout829 _04578_ vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08811_ net602 _05150_ _05116_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_42_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09770__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09791_ _04947_ _06130_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__xnor2_1
Xhold1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[4\] net892 vssd1
+ vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__and3_1
Xhold1027 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[24\] vssd1 vssd1 vccd1 vccd1
+ net2643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2665 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_77_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09522__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08673_ net1073 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[7\] net907 vssd1
+ vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__and3_1
XANTENNA__08876__A2 _04771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08628__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12358__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10667__A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1083_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A _07962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10435__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09225_ net1150 net619 net593 net600 vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout606_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1250_A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_86_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09156_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[16\] net930
+ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07976__A team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11396__B1 _07699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08107_ _04503_ net1161 team_01_WB.instance_to_wrap.cpu.f0.state\[7\] _04577_ vssd1
+ vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__a31o_1
X_09087_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[13\] net926 vssd1
+ vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__and3_1
XANTENNA__12093__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08800__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13137__A1 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08038_ net1661 net568 net346 team_01_WB.instance_to_wrap.cpu.f0.i\[17\] vssd1 vssd1
+ vccd1 vccd1 _03553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold850 _02085_ vssd1 vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold861 _02001_ vssd1 vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[11\] vssd1 vssd1 vccd1 vccd1 net2488
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11010__B net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold883 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold894 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ _06339_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__inv_2
X_09989_ _06325_ _06326_ _06327_ _06328_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__or4_1
XFILLER_0_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10371__A1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1550 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[27\] vssd1 vssd1 vccd1 vccd1
+ net3166 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09513__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1561 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3177 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1572 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3188 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09134__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ net2705 net298 net478 vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1583 team_01_WB.instance_to_wrap.cpu.K0.code\[5\] vssd1 vssd1 vccd1 vccd1 net3199
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1594 team_01_WB.instance_to_wrap.cpu.K0.code\[3\] vssd1 vssd1 vccd1 vccd1 net3210
+ sky130_fd_sc_hd__dlygate4sd3_1
X_10902_ _07003_ _07009_ net519 vssd1 vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__mux2_1
X_11882_ net3025 net283 net485 vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__mux2_1
XANTENNA__11871__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14670_ net1377 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__inv_2
XANTENNA__12776__B _07231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08973__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10833_ _06220_ _07172_ vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__or2_2
XANTENNA__11680__B net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13621_ net187 _04059_ _04060_ net728 vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_120_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12268__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08619__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16340_ clknet_leaf_76_wb_clk_i net2462 _00323_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11623__A1 _07566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13552_ net197 net193 _07816_ _07861_ net643 vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__o2111a_1
X_10764_ net512 net510 _06811_ net511 net538 net544 vssd1 vssd1 vccd1 vccd1 _07104_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_66_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17252__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10977__A3 _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12503_ net2515 net237 net407 vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16271_ clknet_leaf_113_wb_clk_i net1167 _00259_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
X_13483_ _03850_ _03851_ _03943_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10695_ _06902_ _07030_ _07032_ _07034_ _07026_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__o41a_1
X_18010_ net1510 vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_hd__buf_2
XANTENNA__11900__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12434_ net3192 net244 net415 vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__mux2_1
X_15222_ net1200 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__inv_2
XANTENNA__13376__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_81_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15153_ net1291 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__inv_2
X_12365_ net2176 net275 net424 vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13128__A1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14104_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[53\] _04236_ _04244_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[101\]
+ _04390_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__a221o_1
X_11316_ team_01_WB.instance_to_wrap.cpu.f0.state\[8\] _07651_ vssd1 vssd1 vccd1 vccd1
+ _07653_ sky130_fd_sc_hd__or2_1
X_15084_ net1209 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12296_ net2861 net213 net433 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14035_ _04320_ _04321_ _04322_ _04324_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__or4_1
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11247_ _06934_ _07524_ _07583_ vssd1 vssd1 vccd1 vccd1 _07587_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_107_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09752__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09606__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11178_ _07275_ _07515_ _07517_ _07514_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08510__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ _06255_ _06410_ _06441_ _06468_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__a211oi_4
X_15986_ net1384 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__inv_2
X_17725_ clknet_leaf_109_wb_clk_i net871 _01666_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14937_ net1304 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
XANTENNA__09044__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17656_ clknet_leaf_90_wb_clk_i _03341_ _01597_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14868_ net1263 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16607_ clknet_leaf_7_wb_clk_i _02294_ _00590_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13819_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\] net834 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[12\] sky130_fd_sc_hd__and2_1
X_17587_ clknet_leaf_79_wb_clk_i _03274_ _01546_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12178__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14799_ net1214 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13603__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16538_ clknet_leaf_109_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[4\]
+ _00521_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11614__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16469_ clknet_leaf_84_wb_clk_i _02223_ _00452_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11090__A2 _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11810__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09010_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[9\] net911 vssd1
+ vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_94_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold102 _02045_ vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold113 _02005_ vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold124 net111 vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold135 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[4\] vssd1 vssd1 vccd1 vccd1 net1751
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09991__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold146 team_01_WB.instance_to_wrap.a1.ADR_I\[17\] vssd1 vssd1 vccd1 vccd1 net1762
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 net1773
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _02055_ vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ net557 _05264_ net378 vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold179 team_01_WB.instance_to_wrap.a1.ADR_I\[9\] vssd1 vssd1 vccd1 vccd1 net1795
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12641__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout604 _04151_ vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_4
Xfanout615 _07635_ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__clkbuf_4
Xfanout626 net627 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__buf_4
XANTENNA__09743__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09843_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[13\] net802 net784 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__a22o_1
Xfanout637 net638 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__buf_2
XANTENNA__08420__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout648 _04825_ vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout659 net660 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17125__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09774_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[15\] net799 net786 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__a22o_1
XANTENNA__14095__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[5\] net674 _05045_ _05049_
+ _05051_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_59_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08849__A2 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout556_A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1298_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[10\] net680 _04975_
+ _04977_ _04980_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11853__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09889__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17275__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12088__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08587_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[15\] net903
+ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout723_A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10408__A2 _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12802__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09208_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[17\] net897
+ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10480_ _06811_ _06813_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__nor2_1
XANTENNA__09026__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09139_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[14\] net908
+ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08314__B net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ net2765 net300 net452 vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__mux2_1
XANTENNA__09982__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17895__1598 vssd1 vssd1 vccd1 vccd1 net1598 _17895__1598/LO sky130_fd_sc_hd__conb_1
XANTENNA__09129__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11101_ _07161_ _07440_ _07276_ vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__a21o_1
X_12081_ net2617 net284 net462 vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__mux2_1
XANTENNA__12551__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold680 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[28\] vssd1 vssd1 vccd1 vccd1
+ net2307 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08968__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032_ _05417_ net342 vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13530__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08330__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15840_ net1370 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_139_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ net1320 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ net3092 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[111\] net862 vssd1 vssd1
+ vccd1 vccd1 _02142_ sky130_fd_sc_hd__mux2_1
XANTENNA__13294__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1380 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1
+ net2996 sky130_fd_sc_hd__dlygate4sd3_1
X_17510_ clknet_leaf_41_wb_clk_i _03197_ _01493_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14722_ net1316 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__inv_2
Xhold1391 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3007 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_103_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11934_ net2041 net208 net475 vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17441_ clknet_leaf_43_wb_clk_i _03128_ _01424_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14653_ net1241 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__inv_2
X_11865_ net3174 net248 net485 vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16642__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17768__CLK clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_107_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13597__A1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13604_ _03908_ _03900_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__and2b_1
X_17372_ clknet_leaf_37_wb_clk_i _03059_ _01355_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10100__A _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10816_ net510 net509 _06065_ net507 net548 net537 vssd1 vssd1 vccd1 vccd1 _07156_
+ sky130_fd_sc_hd__mux4_2
X_14584_ net1384 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__inv_2
X_11796_ net2836 net213 net491 vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09265__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16323_ clknet_leaf_75_wb_clk_i net1674 _00306_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13535_ net725 _07600_ net980 vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__a21oi_1
X_10747_ _06934_ _07065_ _07079_ _07086_ vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__a211o_1
XANTENNA__11630__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_47 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16254_ clknet_leaf_95_wb_clk_i net1713 _00242_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
X_10678_ _06963_ _06973_ _07016_ _06934_ _06997_ vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__a221o_1
X_13466_ _05655_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 _03927_ sky130_fd_sc_hd__and2b_1
XANTENNA__14010__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10754__B _05996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15205_ net1205 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12417_ net1843 net296 net421 vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16185_ clknet_leaf_112_wb_clk_i _01945_ _00173_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13397_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] _05530_ vssd1 vssd1
+ vccd1 vccd1 _03858_ sky130_fd_sc_hd__or2_1
XANTENNA__08776__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09973__B1 _06311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15136_ net1242 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__inv_2
XANTENNA__08776__B2 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12348_ net2316 net304 net427 vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15338__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ net2454 net227 net437 vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__mux2_1
XANTENNA__12461__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15067_ net1180 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__inv_2
XANTENNA__14242__A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09725__B1 _06063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ _04295_ _04300_ _04305_ _04308_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__or4_2
XANTENNA__11532__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16172__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17298__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15969_ net1334 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10099__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11805__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08510_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[18\] net893 vssd1
+ vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__and3_1
X_17708_ clknet_leaf_101_wb_clk_i _03392_ _01649_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[29\]
+ sky130_fd_sc_hd__dfrtp_2
X_09490_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[30\] net700 _05829_ net706
+ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08700__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[23\] net910
+ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17639_ clknet_leaf_111_wb_clk_i _03324_ _01580_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09502__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08372_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__nor2_2
XANTENNA__15801__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09110__D1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12636__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14001__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout304_A _07912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10023__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1046_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12371__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13512__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 _03566_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_8
Xfanout412 _03563_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__buf_4
XANTENNA__16515__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09716__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11495__B net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout423 _07966_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_8
Xfanout434 _07964_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 _07959_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout673_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout456 _07956_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_4
X_09826_ net1134 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[13\] net959
+ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout467 net470 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_35_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout478 _07950_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout489 _07947_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_8
XFILLER_0_96_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout840_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\] net764 net621 vssd1
+ vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13276__B1 _07650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout938_A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11715__S net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[5\] net909 vssd1
+ vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09688_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[22\] net746 _06004_ _06008_
+ _06009_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_16_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08639_ net1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[10\] net896
+ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08309__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11016__A _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10558__C net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11650_ _07856_ _07857_ net611 vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__mux2_4
XANTENNA__09247__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10601_ _06939_ _06940_ vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11581_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] _07797_ vssd1 vssd1 vccd1
+ vccd1 _07798_ sky130_fd_sc_hd__and2_1
XANTENNA__12546__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10855__A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10532_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[31\] net655 net649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__a22o_1
X_13320_ net565 _07706_ _07731_ net829 vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__a31o_1
XFILLER_0_52_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10463_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[26\] net799 net762 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__a22o_1
X_13251_ _07686_ _07702_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__nor2_1
XANTENNA__13200__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12202_ net2527 net273 net445 vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13182_ net1164 team_01_WB.instance_to_wrap.a1.prev_BUSY_O net835 vssd1 vssd1 vccd1
+ vccd1 _03738_ sky130_fd_sc_hd__and3b_2
X_10394_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[16\] net824 _06732_ _06733_
+ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__a211o_1
XANTENNA_input67_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12133_ net2935 net205 net451 vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12281__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15158__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17990_ net1490 vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__buf_2
XANTENNA__16195__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13503__A1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09156__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ net2713 net247 net461 vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__mux2_1
X_16941_ clknet_leaf_140_wb_clk_i _02628_ _00924_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11015_ _05594_ net508 vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_109_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16872_ clknet_leaf_30_wb_clk_i _02559_ _00855_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout990 _04491_ vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__clkbuf_2
X_15823_ net1322 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11625__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15754_ net1400 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__inv_2
X_12966_ net1161 team_01_WB.instance_to_wrap.cpu.f0.state\[3\] vssd1 vssd1 vccd1 vccd1
+ _03718_ sky130_fd_sc_hd__nand2_1
XANTENNA__09486__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ net1319 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11917_ net2451 net282 net479 vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15685_ net1207 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__inv_2
X_12897_ net361 _03672_ net1029 vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_64_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17424_ clknet_leaf_126_wb_clk_i _03111_ _01407_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14636_ net1216 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ net3214 net254 net489 vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__mux2_1
XANTENNA__09238__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17355_ clknet_leaf_3_wb_clk_i _03042_ _01338_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12242__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14567_ net1338 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11779_ net2655 net227 net496 vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16306_ clknet_leaf_61_wb_clk_i _02060_ _00289_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[29\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13518_ net722 _07566_ net1066 vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__o21a_1
X_17286_ clknet_leaf_40_wb_clk_i _02973_ _01269_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14498_ net1383 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16237_ clknet_leaf_105_wb_clk_i net1888 _00225_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_1
X_13449_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _04946_ _03902_ vssd1
+ vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_77_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_75_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10005__B1 _04684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16538__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16168_ clknet_leaf_102_wb_clk_i net3148 _00156_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09410__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10556__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11596__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15119_ net1216 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15068__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12191__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08990_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[8\] net923 vssd1
+ vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__and3_1
X_16099_ clknet_leaf_83_wb_clk_i _01874_ _00087_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10859__A2 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09611_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[24\] net789 net754 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09542_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[28\] net954
+ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_1590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09477__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09473_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[30\] net926 vssd1
+ vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_138_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout254_A _07904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17894__1597 vssd1 vssd1 vccd1 vccd1 net1597 _17894__1597/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_138_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08424_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[23\] net931
+ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_138_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[30\] net818 net760 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[30\]
+ _04694_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12366__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13430__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17313__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1163_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10244__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08286_ net1156 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__or3b_2
XANTENNA__10795__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1330_A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07984__A team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13733__A1 team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13733__B2 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout790_A _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17463__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09401__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout888_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11744__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1207 net1208 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__buf_4
Xfanout1218 net1236 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__buf_2
XANTENNA__13497__B1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout220 net221 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_2
Xfanout1229 net1231 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__buf_4
Xfanout231 net234 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_2
Xfanout242 _07870_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_1
Xfanout253 _07904_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_2
Xfanout264 net266 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_2
Xfanout275 net277 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_2
Xfanout286 _07908_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_2
X_09809_ _06141_ _06142_ _06143_ _06148_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__or4_1
Xfanout297 _07926_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12820_ net366 _03641_ _03642_ net1057 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__a32o_1
XFILLER_0_119_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12751_ net1025 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[25\] vssd1 vssd1 vccd1
+ vccd1 _03595_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11702_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] _07803_ vssd1 vssd1
+ vccd1 vccd1 _07899_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15470_ net1282 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__inv_2
X_12682_ net3010 net310 net390 vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08981__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ net1360 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[25\] net715 net616 vssd1 vssd1
+ vccd1 vccd1 _07844_ sky130_fd_sc_hd__o21a_1
XANTENNA__12276__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17140_ clknet_leaf_128_wb_clk_i _02827_ _01123_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14352_ net1363 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__inv_2
X_11564_ team_01_WB.instance_to_wrap.cpu.K0.count\[1\] team_01_WB.instance_to_wrap.cpu.K0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__nand2_1
XFILLER_0_52_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13303_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] net610 _07707_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__a31o_1
X_17071_ clknet_leaf_143_wb_clk_i _02758_ _01054_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10515_ _06847_ _06848_ _06853_ _06854_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__or4_4
XFILLER_0_68_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11495_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[15\] net580 vssd1 vssd1 vccd1
+ vccd1 _07775_ sky130_fd_sc_hd__nand2_1
X_14283_ net1374 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__inv_2
XANTENNA__09928__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16022_ net1375 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__inv_2
X_10446_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[26\] net968
+ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__and3b_1
X_13234_ net2367 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1
+ vccd1 vccd1 _01916_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10538__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10377_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[16\] net959
+ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__and3_1
X_13165_ net1820 net843 net840 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[11\] vssd1
+ vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a22o_1
X_17928__1616 vssd1 vssd1 vccd1 vccd1 net1616 _17928__1616/LO sky130_fd_sc_hd__conb_1
X_12116_ net1884 net280 net456 vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__mux2_1
X_17973_ net1473 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
X_13096_ net50 net39 net64 net61 vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__or4_1
XFILLER_0_137_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16924_ clknet_leaf_37_wb_clk_i _02611_ _00907_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12047_ net1882 net253 net463 vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16855_ clknet_leaf_137_wb_clk_i _02542_ _00838_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16980__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15806_ net1352 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_122_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_66_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16786_ clknet_leaf_129_wb_clk_i _02473_ _00769_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13998_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\]
+ _04237_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_66_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15737_ net1261 vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__inv_2
XANTENNA__09052__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[7\] net1036 vssd1 vssd1 vccd1
+ vccd1 _03709_ sky130_fd_sc_hd__nor2_1
XANTENNA__16210__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10198__C net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17336__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15668_ net1267 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__inv_2
XANTENNA__08891__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17407_ clknet_leaf_7_wb_clk_i _03094_ _01390_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14619_ net1375 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__inv_2
XANTENNA__12186__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15599_ net1217 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08140_ _04606_ _04607_ _04608_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17338_ clknet_leaf_60_wb_clk_i _03025_ _01321_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12766__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11423__C1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10777__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17486__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08071_ _04515_ _04523_ _04537_ _04546_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__or4_2
X_17269_ clknet_leaf_125_wb_clk_i _02956_ _01252_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09495__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09919__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09395__A1 _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13191__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08412__B net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[8\] net923 vssd1
+ vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold17 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[80\] vssd1 vssd1 vccd1 vccd1 net1633
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold28 _03529_ vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold39 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[7\] vssd1 vssd1 vccd1 vccd1 net1655
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout469_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11065__A2_N net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09525_ _05855_ _05860_ _05864_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__nor3_1
XFILLER_0_79_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1280_A net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1378_A net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_26_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09456_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[29\] net699 net692 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[29\]
+ _05786_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_26_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09870__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08407_ _04738_ _04745_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__and2b_1
XFILLER_0_137_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12096__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10609__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout803_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] net712 net594 vssd1 vssd1
+ vccd1 vccd1 _05727_ sky130_fd_sc_hd__a21o_1
XANTENNA__13403__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10217__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12757__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08338_ net1134 net959 vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_95_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08269_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[12\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\]
+ net1038 vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10300_ net505 _06638_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__or2_1
X_11280_ _07054_ _07497_ _07614_ _06963_ _07619_ vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__a221o_1
X_10231_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[9\] net745 net741 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10162_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] net626 vssd1 vssd1 vccd1
+ vccd1 _06502_ sky130_fd_sc_hd__nand2_2
XFILLER_0_98_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09137__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1004 net1009 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1015 net1016 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__buf_2
XFILLER_0_105_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1026 net1029 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_2
Xfanout1037 net1038 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__clkbuf_4
X_10093_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[7\] net812 net779 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[7\]
+ _06411_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__a221o_1
X_14970_ net1192 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__inv_2
Xfanout1048 net1049 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_2
Xfanout1059 team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1 vccd1
+ net1059 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13921_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\]
+ _04212_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__and3_1
XANTENNA__08976__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16233__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16640_ clknet_leaf_33_wb_clk_i _02327_ _00623_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08361__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13852_ net1166 net1060 net1721 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[13\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_18_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12803_ net1795 net641 net608 _03630_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a22o_1
X_16571_ clknet_leaf_54_wb_clk_i _02258_ _00554_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_13783_ _04162_ _01835_ _04166_ _04159_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__o211a_1
X_10995_ net563 net338 _07334_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11903__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15522_ net1312 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__inv_2
X_12734_ net2361 net642 _03582_ net606 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09861__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15453_ net1262 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__inv_2
X_12665_ net3002 net243 net387 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14404_ net1332 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11616_ net616 _07830_ _07829_ vssd1 vssd1 vccd1 vccd1 _07831_ sky130_fd_sc_hd__o21ai_4
X_15384_ net1183 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12596_ net2039 net274 net397 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__mux2_1
XANTENNA__09613__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17123_ clknet_leaf_23_wb_clk_i _02810_ _01106_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14335_ net1377 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__inv_2
X_11547_ net2511 net1160 vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17054_ clknet_leaf_44_wb_clk_i _02741_ _01037_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold509 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14266_ net1317 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11478_ net367 _07766_ net3100 net874 vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08513__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16005_ net1353 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__inv_2
XANTENNA__13173__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13217_ net566 _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10429_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[27\] net783 _06755_ _06759_
+ _06762_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_1404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14197_ net1734 _04462_ net1410 vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11184__A1 _07014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17893__1596 vssd1 vssd1 vccd1 vccd1 net1596 _17893__1596/LO sky130_fd_sc_hd__conb_1
XANTENNA__12920__A2 _03688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13148_ net1698 net845 net839 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[28\] vssd1
+ vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09047__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15346__A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13079_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\] net3113 net863 vssd1 vssd1
+ vccd1 vccd1 _02046_ sky130_fd_sc_hd__mux2_1
X_17956_ net1456 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
Xhold1209 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08886__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09344__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16907_ clknet_leaf_3_wb_clk_i _02594_ _00890_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_17887_ net107 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08352__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16838_ clknet_leaf_40_wb_clk_i _02525_ _00821_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16726__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16769_ clknet_leaf_41_wb_clk_i _02456_ _00752_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_124_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11813__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09310_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[22\] net665 _05627_
+ _05629_ _05641_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_130_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09241_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[21\] net672 net649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09510__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16876__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_90_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09172_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[16\] net906
+ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ _04480_ team_01_WB.instance_to_wrap.cpu.f0.num\[14\] team_01_WB.instance_to_wrap.cpu.f0.num\[13\]
+ _04481_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_86_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12644__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08812__B1 _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout217_A _07835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08054_ team_01_WB.instance_to_wrap.cpu.K0.code\[7\] team_01_WB.instance_to_wrap.cpu.K0.code\[6\]
+ team_01_WB.instance_to_wrap.cpu.K0.code\[4\] team_01_WB.instance_to_wrap.cpu.K0.code\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__or4b_2
XANTENNA__08423__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_133_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13164__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11175__A1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1126_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10367__A1_N net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16256__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08591__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _05292_ _05293_ _05294_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__or4_1
XANTENNA__17501__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08796__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08879__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[2\] net921 vssd1
+ vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout753_A _04678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10150__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout920_A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09508_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[29\] net973
+ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10780_ net515 _07105_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17927__1615 vssd1 vssd1 vccd1 vccd1 net1615 _17927__1615/LO sky130_fd_sc_hd__conb_1
XANTENNA__09843__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09439_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\] net704 _05774_ _05778_
+ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__o22a_4
XFILLER_0_94_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08317__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12450_ net2499 net294 net418 vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__mux2_1
X_11401_ _07696_ _07714_ team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1
+ vccd1 _07724_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12381_ net2136 net302 net425 vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__mux2_1
XANTENNA__12554__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14120_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[86\] _04251_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[118\]
+ _04397_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11332_ _07664_ net1758 _07655_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__mux2_1
XANTENNA__08333__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10582__B _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14054__B _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14051_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[75\] _04235_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[123\]
+ _04339_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__a221o_1
X_11263_ net529 _07106_ vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_123_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13002_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[84\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[92\]
+ net856 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__mux2_1
X_10214_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[8\] net747 _06537_ _06541_
+ _06543_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__a2111o_1
X_11194_ _07058_ _07080_ net514 vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__mux2_1
XANTENNA__08031__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_105_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17181__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17810_ clknet_leaf_85_wb_clk_i _03486_ _01750_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[80\]
+ sky130_fd_sc_hd__dfrtp_1
X_10145_ _06481_ _06482_ _06483_ _06484_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17741_ clknet_leaf_77_wb_clk_i net2759 _01681_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09164__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16749__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14953_ net1228 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__inv_2
X_10076_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[7\] net959 vssd1
+ vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__and3_1
X_13904_ _04204_ net571 _04203_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__and3b_1
XANTENNA__10677__B1 _06921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17672_ clknet_leaf_119_wb_clk_i _03357_ _01613_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10103__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14884_ net1237 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
XANTENNA__10141__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16623_ clknet_leaf_144_wb_clk_i _02310_ _00606_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13835_ net1697 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[28\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_98_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13414__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16554_ clknet_leaf_116_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[20\]
+ _00537_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13766_ _04154_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ _06438_ net373 net550 vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__mux2_1
XANTENNA__08508__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09834__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15505_ net1288 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__inv_2
X_12717_ net2808 net319 net386 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16485_ clknet_leaf_95_wb_clk_i _02239_ _00468_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13697_ _04110_ _04111_ _04119_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[15\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_128_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15436_ net1219 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__inv_2
X_12648_ net2781 net296 net394 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_84_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_81_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15367_ net1325 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12464__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12579_ net2399 net304 net400 vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14245__A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17106_ clknet_leaf_130_wb_clk_i _02793_ _01089_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14318_ net1347 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08270__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_18086_ net636 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
Xhold306 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15298_ net1264 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__inv_2
Xhold317 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[56\] vssd1 vssd1 vccd1 vccd1
+ net1933 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 _01987_ vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[9\] vssd1 vssd1 vccd1 vccd1 net1955
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13146__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17037_ clknet_leaf_2_wb_clk_i _02724_ _01020_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14249_ net1354 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11157__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout808 net810 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__buf_8
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout819 _04632_ vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_8
X_08810_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] net702 _05133_ _05149_
+ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__o22a_4
XANTENNA__11808__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ _04969_ _05378_ _05492_ net561 vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__a31o_1
Xhold1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10380__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1017 team_01_WB.instance_to_wrap.cpu.K0.count\[1\] vssd1 vssd1 vccd1 vccd1 net2633
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[4\] net909 vssd1
+ vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__and3_1
XANTENNA__17674__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12657__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17939_ net1439 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
Xhold1028 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09505__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1390 net1391 vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__buf_4
XANTENNA__15804__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08672_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[7\] net934 vssd1
+ vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08730__C1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12639__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10667__B _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08418__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout334_A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10840__A0 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1076_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09224_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] net702 _05561_ _05563_
+ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__o22a_4
XFILLER_0_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14031__B1 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09155_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] net619 net593 vssd1 vssd1
+ vccd1 vccd1 _05495_ sky130_fd_sc_hd__a21o_1
XANTENNA__12374__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout501_A _07795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1243_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08106_ _04511_ _04575_ _04576_ net1036 vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__o31a_1
XFILLER_0_27_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09086_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[13\] net910
+ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13137__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08037_ net1736 net567 net346 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1
+ vccd1 vccd1 _03554_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1410_A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold840 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[32\] vssd1 vssd1 vccd1 vccd1
+ net2456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold851 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold862 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13542__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold873 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold884 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[6\] vssd1 vssd1 vccd1 vccd1
+ net2511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08564__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11718__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[2\] net796 _04654_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_129_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08939_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[6\] net880 vssd1
+ vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__and3_1
XANTENNA__12648__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17989__1489 vssd1 vssd1 vccd1 vccd1 _17989__1489/HI net1489 sky130_fd_sc_hd__conb_1
Xhold1540 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net3156 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10659__A0 _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1551 _03441_ vssd1 vssd1 vccd1 vccd1 net3167 sky130_fd_sc_hd__dlygate4sd3_1
X_11950_ net1880 net282 net475 vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__mux2_1
Xhold1562 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3178 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10123__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1573 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1584 team_01_WB.instance_to_wrap.cpu.K0.code\[2\] vssd1 vssd1 vccd1 vccd1 net3200
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1595 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net3211 sky130_fd_sc_hd__dlygate4sd3_1
X_10901_ net523 _07240_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__or2_1
X_11881_ net1966 net253 net484 vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__mux2_1
XANTENNA__12549__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13620_ net199 net195 _07804_ _07903_ net645 vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_120_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10832_ _06469_ _06472_ _06597_ _06603_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_120_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08328__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13551_ _03932_ _04001_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__xnor2_1
X_17892__1595 vssd1 vssd1 vccd1 vccd1 net1595 _17892__1595/LO sky130_fd_sc_hd__conb_1
X_10763_ _06958_ _07099_ _07102_ _07098_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12820__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12502_ net2937 net240 net407 vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16270_ clknet_leaf_4_wb_clk_i _02030_ _00258_ vssd1 vssd1 vccd1 vccd1 team_01_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10831__B1 _07170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14022__B1 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _05679_ _05705_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\]
+ _03941_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__a221o_1
X_10694_ _06906_ _07033_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15221_ net1223 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__inv_2
XANTENNA__13376__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12433_ net2632 net202 net415 vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__mux2_1
XANTENNA__12284__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16421__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15152_ net1272 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12364_ net2154 net211 net426 vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_105_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14103_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[45\] _04246_ _04251_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[85\]
+ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13128__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11315_ team_01_WB.instance_to_wrap.cpu.f0.state\[8\] _07651_ vssd1 vssd1 vccd1 vccd1
+ _07652_ sky130_fd_sc_hd__nor2_2
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15083_ net1295 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12295_ net2306 net219 net433 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__mux2_1
X_14034_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[26\] _04243_ _04254_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[98\]
+ _04323_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__a221o_1
XANTENNA__13533__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11246_ net555 _07528_ _07582_ _07345_ _07585_ vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12887__A1 _03665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17697__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08555__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13409__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11177_ net531 _07445_ _07516_ net330 vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10362__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10128_ net373 _06467_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__and2_1
X_15985_ net1333 vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10059_ net550 _06398_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__or2_1
XANTENNA__15624__A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17724_ clknet_leaf_109_wb_clk_i _00006_ _01665_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_14936_ net1183 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10114__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14867_ net1278 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
XANTENNA__11464__A2_N net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17655_ clknet_leaf_90_wb_clk_i _03340_ _01596_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12459__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16606_ clknet_leaf_48_wb_clk_i _02293_ _00589_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13818_ net1798 net834 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[11\]
+ sky130_fd_sc_hd__and2_1
X_17586_ clknet_leaf_79_wb_clk_i _03273_ _01545_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09268__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14798_ net1283 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__inv_2
XANTENNA__09807__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16537_ clknet_leaf_90_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[3\]
+ _00520_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12811__A1 _07323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09060__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11614__A2 _07056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13749_ _04115_ team_01_WB.instance_to_wrap.cpu.c0.next_count\[16\] _04138_ team_01_WB.instance_to_wrap.cpu.c0.next_count\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_atmax sky130_fd_sc_hd__and4b_1
XFILLER_0_50_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16468_ clknet_leaf_136_wb_clk_i _02222_ _00451_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14013__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11599__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15419_ net1181 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__inv_2
XANTENNA__12194__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16399_ clknet_leaf_67_wb_clk_i net1905 _00382_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16914__CLK clknet_leaf_132_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold103 net95 vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13119__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold114 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[12\] vssd1 vssd1 vccd1 vccd1
+ net1730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold125 _01978_ vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
X_18069_ net1569 vssd1 vssd1 vccd1 vccd1 la_data_out[111] sky130_fd_sc_hd__buf_2
Xhold136 _01970_ vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12922__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold147 _02015_ vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold158 team_01_WB.instance_to_wrap.cpu.f0.write_data\[7\] vssd1 vssd1 vccd1 vccd1
+ net1774 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _06250_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold169 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12878__A1 _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout605 _04151_ vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__dlymetal6s2s_1
X_17926__1614 vssd1 vssd1 vccd1 vccd1 net1614 _17926__1614/LO sky130_fd_sc_hd__conb_1
Xfanout616 _07635_ vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_8
X_09842_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[13\] net785 net740 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[13\]
+ _06181_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout627 _04627_ vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_8
Xfanout638 net179 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout649 _04823_ vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__buf_6
XANTENNA__08420__B net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10353__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[15\] net792 net752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[15\]
+ _06112_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_52_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[5\] net700 net669 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10105__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09532__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08655_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[10\] net671 _04989_ _04993_
+ _04994_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_94_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12369__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout451_A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1193_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout549_A _05151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09259__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08586_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[15\] net937 vssd1
+ vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12802__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16444__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07987__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14004__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09207_ net1075 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[17\] net905
+ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09138_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[14\] net902
+ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16594__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09431__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09069_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[12\] net692 _05384_ _05395_
+ _05403_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_130_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11100_ _06921_ _07160_ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12080_ net2925 net252 net460 vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__mux2_1
XANTENNA__12869__A1 _06881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[20\] vssd1 vssd1 vccd1 vccd1 net2308
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ _07369_ _07370_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13530__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15770_ net1316 vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[104\] net2534 net863 vssd1 vssd1
+ vccd1 vccd1 _02143_ sky130_fd_sc_hd__mux2_1
XANTENNA__13294__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1370 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[82\] vssd1 vssd1 vccd1 vccd1
+ net2986 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14721_ net1316 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__inv_2
Xhold1381 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11933_ net2878 net275 net477 vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__mux2_1
XANTENNA__12279__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1392 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3008 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_103_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17440_ clknet_leaf_33_wb_clk_i _03127_ _01423_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14652_ net1254 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__inv_2
X_11864_ net1930 net215 net484 vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13603_ net981 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] _04044_ _04045_
+ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a22o_1
X_17371_ clknet_leaf_17_wb_clk_i _03058_ _01354_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10815_ _06106_ _06744_ _06747_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__nand3_1
XANTENNA__13597__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14583_ net1339 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11795_ net2596 net216 net491 vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__mux2_1
XANTENNA__11911__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16322_ clknet_leaf_61_wb_clk_i _02076_ _00305_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[45\]
+ sky130_fd_sc_hd__dfstp_1
X_13534_ net185 _03986_ _03987_ net725 vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__a211o_1
XFILLER_0_138_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10746_ net523 _07082_ _07083_ _05263_ _07085_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16253_ clknet_leaf_84_wb_clk_i _02013_ _00241_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_125_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13465_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] _04842_ vssd1 vssd1
+ vccd1 vccd1 _03926_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10677_ net554 _06858_ _06921_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_11_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15204_ net1237 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__inv_2
X_12416_ net3077 net298 net421 vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16184_ clknet_leaf_107_wb_clk_i _01944_ _00172_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13396_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] _05530_ vssd1 vssd1
+ vccd1 vccd1 _03857_ sky130_fd_sc_hd__and2_1
XANTENNA__09422__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09973__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15135_ net1254 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12347_ net2601 net286 net430 vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__mux2_1
XANTENNA__15619__A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13506__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15066_ net1191 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__inv_2
X_12278_ net2973 net288 net438 vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08521__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14017_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[49\] _04236_ _04290_ _04307_
+ _04152_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09725__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ _05965_ _07568_ _05934_ vssd1 vssd1 vccd1 vccd1 _07569_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11532__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09055__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09489__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13285__A1 _04621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15968_ net1336 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__inv_2
XANTENNA__08894__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18059__1559 vssd1 vssd1 vccd1 vccd1 _18059__1559/HI net1559 sky130_fd_sc_hd__conb_1
XFILLER_0_91_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17707_ clknet_leaf_103_wb_clk_i _03391_ _01648_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[28\]
+ sky130_fd_sc_hd__dfrtp_4
X_14919_ net1328 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
XANTENNA__12189__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15899_ net1397 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__inv_2
XANTENNA__10498__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08697__D1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16467__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08440_ net1081 net909 vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__and2_2
XFILLER_0_8_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08700__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17638_ clknet_leaf_113_wb_clk_i _03323_ _01579_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08371_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__or4bb_4
X_17569_ clknet_leaf_60_wb_clk_i _03256_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11821__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17988__1488 vssd1 vssd1 vccd1 vccd1 _17988__1488/HI net1488 sky130_fd_sc_hd__conb_1
XFILLER_0_5_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09413__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08767__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15529__A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12652__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1039_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08431__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_A _07795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 _03566_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_4
Xfanout413 _03563_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17891__1594 vssd1 vssd1 vccd1 vccd1 net1594 _17891__1594/LO sky130_fd_sc_hd__conb_1
Xfanout424 _07966_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1206_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 _07963_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout446 _07959_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_4
XANTENNA__11523__B2 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17242__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _06134_ _06164_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__or2_1
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 _07956_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_6
Xfanout468 net470 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout479 _07949_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_6
XANTENNA_fanout666_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ net770 _06089_ _06093_ _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__nor4_1
X_08707_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[5\] net916 vssd1
+ vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__and3_1
XANTENNA__12099__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09687_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[22\] net782 net760 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout833_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17392__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08638_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[10\] net901
+ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11016__B net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08569_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[19\] net878 vssd1
+ vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10600_ net546 net340 vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12787__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11580_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\]
+ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1 _07797_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_119_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10855__B net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10531_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[31\] net694 net687 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13250_ net1939 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1
+ vccd1 vccd1 _01900_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10462_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[26\] net792 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__a22o_1
XANTENNA__09404__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12201_ net1861 net245 net443 vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__mux2_1
XANTENNA__15439__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13181_ team_01_WB.instance_to_wrap.a1.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1
+ _03737_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12562__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10393_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[16\] net804 net755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12132_ net2604 net275 net451 vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10970__C1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13503__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12063_ net2528 net214 net461 vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__mux2_1
X_16940_ clknet_leaf_133_wb_clk_i _02627_ _00923_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10317__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11514__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11496__A1_N net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11014_ _05595_ net508 vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_109_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16871_ clknet_leaf_123_wb_clk_i _02558_ _00854_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout980 net981 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__buf_2
XANTENNA__11906__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15822_ net1317 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout991 net993 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__buf_2
XANTENNA__17735__CLK clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13267__B2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09172__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17910__1602 vssd1 vssd1 vccd1 vccd1 net1602 _17910__1602/LO sky130_fd_sc_hd__conb_1
X_15753_ net1400 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__inv_2
X_12965_ net2015 net873 net360 _03717_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a22o_1
XANTENNA__09603__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15902__A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11916_ net2485 net304 net481 vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ net1318 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__inv_2
X_15684_ net1238 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _04837_ net577 vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ net1297 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__inv_2
XANTENNA__17885__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17423_ clknet_leaf_143_wb_clk_i _03110_ _01406_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ net2664 net227 net489 vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14518__A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925__1613 vssd1 vssd1 vccd1 vccd1 net1613 _17925__1613/LO sky130_fd_sc_hd__conb_1
X_14566_ net1337 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__inv_2
X_17354_ clknet_leaf_11_wb_clk_i _03041_ _01337_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11778_ net1902 net290 net497 vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08516__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16305_ clknet_leaf_59_wb_clk_i _02059_ _00288_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[28\]
+ sky130_fd_sc_hd__dfstp_1
X_13517_ net185 _03972_ _03973_ net725 vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17285_ clknet_leaf_39_wb_clk_i _02972_ _01268_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10729_ _06920_ _06928_ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17115__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13990__A2 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14497_ net1396 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16236_ clknet_leaf_105_wb_clk_i net1704 _00224_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_1
X_13448_ _03904_ _03907_ _03908_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__nand3_1
XFILLER_0_109_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12472__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16167_ clknet_leaf_97_wb_clk_i _01930_ _00155_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13379_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] _05834_ vssd1 vssd1
+ vccd1 vccd1 _03840_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_58_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11753__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15118_ net1284 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__inv_2
XANTENNA__08889__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11596__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17265__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16098_ clknet_leaf_93_wb_clk_i _01873_ _00086_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15049_ net1230 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09174__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10859__A3 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11816__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09610_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[24\] net758 _05936_ _05942_
+ _05945_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_121_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08921__A2 _05258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09082__A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09541_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[28\] net968 vssd1
+ vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11117__A _06921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09472_ net1071 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[30\] net897
+ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_138_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08423_ net1083 net930 vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_138_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12647__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10956__A _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12769__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08354_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[30\] net785 net735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13430__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08426__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11441__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13981__A2 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08285_ _04623_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout414_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13194__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12382__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10691__A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1323_A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08799__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout783_A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1208 net1211 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__buf_4
XANTENNA__13497__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout210 net212 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_2
Xfanout1219 net1227 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__buf_4
Xfanout221 _07831_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_2
Xfanout232 net234 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09165__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout243 _07862_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_2
Xfanout254 _07904_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_2
Xfanout276 net277 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08912__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ _06144_ _06145_ _06146_ _06147_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__or4_1
Xfanout287 net290 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_2
XANTENNA__10180__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout298 net301 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_2
Xclkbuf_4_15__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_104_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13249__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16782__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09739_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[20\] net964
+ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12750_ net1027 net278 vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11701_ net721 _07207_ net615 _07897_ vssd1 vssd1 vccd1 vccd1 _07898_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12681_ net2558 net296 net388 vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__mux2_1
XANTENNA__12557__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17138__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14420_ net1366 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ net716 net278 vssd1 vssd1 vccd1 vccd1 _07843_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08979__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14351_ net1371 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11432__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11563_ net2859 net1168 net34 vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13302_ net1658 net825 _03783_ _03785_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__o22a_1
XANTENNA__10786__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10514_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[31\] net790 net768 _06837_
+ _06842_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__a2111o_1
XANTENNA__16162__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17070_ clknet_leaf_5_wb_clk_i _02757_ _01053_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17288__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14282_ net1375 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__inv_2
X_11494_ net367 _07774_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[16\] net874
+ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_122_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13185__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16021_ net1356 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13233_ net2855 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[17\] vssd1 vssd1
+ vccd1 vccd1 _01917_ sky130_fd_sc_hd__a22o_1
XANTENNA__11697__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12292__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10445_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[26\] net942
+ vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18058__1558 vssd1 vssd1 vccd1 vccd1 _18058__1558/HI net1558 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_72_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09167__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13164_ net1740 net851 net842 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[12\] vssd1
+ vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10376_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[16\] net969
+ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12115_ net2128 net302 net456 vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__mux2_1
X_17972_ net1472 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_104_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13095_ net66 net65 net68 net67 vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__or4_1
XANTENNA__13488__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12046_ net2747 net229 net463 vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__mux2_1
X_16923_ clknet_leaf_53_wb_clk_i _02610_ _00906_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13417__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16854_ clknet_leaf_1_wb_clk_i _02541_ _00837_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10171__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17987__1487 vssd1 vssd1 vccd1 vccd1 _17987__1487/HI net1487 sky130_fd_sc_hd__conb_1
X_15805_ net1323 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13997_ net1777 net604 _04288_ net1169 vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__o211a_1
X_16785_ clknet_leaf_15_wb_clk_i _02472_ _00768_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12948_ net359 _03707_ _03708_ net872 net3268 vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a32o_1
X_15736_ net1177 vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__inv_2
XANTENNA__09864__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13660__A1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09630__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11671__A0 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15667_ net1280 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__inv_2
X_12879_ net2556 net871 net358 _03660_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__a22o_1
XANTENNA__12467__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17406_ clknet_leaf_46_wb_clk_i _03093_ _01389_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14618_ net1361 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__inv_2
X_15598_ net1283 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
XANTENNA__10495__B net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17337_ clknet_leaf_58_wb_clk_i _03024_ _01320_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14549_ net1395 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10777__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08070_ _04537_ _04546_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17268_ clknet_leaf_128_wb_clk_i _02955_ _01251_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13176__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16219_ clknet_leaf_78_wb_clk_i net1900 _00207_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17199_ clknet_leaf_142_wb_clk_i _02886_ _01182_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10529__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12923__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap977 _04631_ vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09508__C net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10934__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08412__C net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08972_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[8\] net892 vssd1
+ vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__and3_1
XANTENNA__09147__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold18 _02119_ vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14140__A2 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold29 team_01_WB.instance_to_wrap.cpu.f0.write_data\[0\] vssd1 vssd1 vccd1 vccd1
+ net1645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08355__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout197_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout364_A _03580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09524_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[29\] net783 _05861_ _05862_
+ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_79_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09855__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09540__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[29\] net695 _05792_
+ _05793_ _05794_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout531_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12377__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1273_A net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08406_ _04741_ _04744_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09386_ _05713_ _05718_ _05725_ net704 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__o32a_4
XANTENNA__13403__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17430__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08337_ net1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[30\] net948
+ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\]
+ net1040 vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13167__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout998_A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08199_ net2568 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[74\] net1043 vssd1 vssd1
+ vccd1 vccd1 _03488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10230_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[9\] net971 vssd1
+ vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08594__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ _06499_ _06500_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__nor2_1
XANTENNA__12840__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1005 net1006 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_7_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1016 net1017 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1027 net1029 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__buf_2
X_17924__1612 vssd1 vssd1 vccd1 vccd1 net1612 _17924__1612/LO sky130_fd_sc_hd__conb_1
Xfanout1038 net1045 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_2
X_10092_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[7\] net802 net756 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__a22o_1
Xfanout1049 net1053 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__buf_2
XFILLER_0_41_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13920_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\] _04142_ _04207_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13851_ net1166 net1060 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[12\] sky130_fd_sc_hd__and3b_1
XFILLER_0_57_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12802_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] net1056 net365 _03629_
+ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13782_ _04162_ _04165_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__nand2_1
X_16570_ clknet_leaf_59_wb_clk_i _02257_ _00553_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10994_ _06399_ _07010_ vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__nand2_1
XANTENNA__11102__C1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13642__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16528__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08992__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12733_ net1054 team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] net639 vssd1 vssd1
+ vccd1 vccd1 _03583_ sky130_fd_sc_hd__o21ba_1
X_15521_ net1246 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09310__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12287__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11653__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15452_ net1175 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__inv_2
X_12664_ net2285 net203 net387 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14403_ net1403 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__inv_2
X_11615_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] _07820_ vssd1 vssd1
+ vccd1 vccd1 _07830_ sky130_fd_sc_hd__xnor2_2
XANTENNA_clkbuf_leaf_74_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15383_ net1198 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__inv_2
XANTENNA__16678__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12595_ net2842 net209 net397 vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__mux2_1
XANTENNA__11956__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17122_ clknet_leaf_32_wb_clk_i _02809_ _01105_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14334_ net1370 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11546_ net2185 net1159 net589 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1
+ vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13158__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17053_ clknet_leaf_49_wb_clk_i _02740_ _01036_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14265_ net1317 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11477_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[24\] net579 vssd1 vssd1 vccd1
+ vccd1 _07766_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_55_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16004_ net1356 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__inv_2
X_13216_ _04505_ team_01_WB.instance_to_wrap.cpu.f0.state\[6\] _07649_ vssd1 vssd1
+ vccd1 vccd1 _03740_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09377__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10428_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[27\] net822 net751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[27\]
+ _06767_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__a221o_1
X_14196_ net1410 _04461_ _04462_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__nor3_1
XFILLER_0_104_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13147_ net1907 net845 net840 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[29\] vssd1
+ vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__a22o_1
X_10359_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[17\] net775 net772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__a22o_1
XANTENNA__10392__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14122__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09625__A _05963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13078_ net2623 net1783 net860 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__mux2_1
X_17955_ net1455 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
XANTENNA__13851__A_N net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17303__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12029_ net2819 net216 net465 vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__mux2_1
X_16906_ clknet_leaf_11_wb_clk_i _02593_ _00889_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_68_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10144__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17886_ net107 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10695__A1 _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16837_ clknet_leaf_39_wb_clk_i _02524_ _00820_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09063__C _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16768_ clknet_leaf_33_wb_clk_i _02455_ _00751_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13633__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17453__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15719_ net1328 vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11644__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12197__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16699_ clknet_leaf_19_wb_clk_i _02386_ _00682_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09240_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[21\] net677 net653 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[21\]
+ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09171_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[16\] net930 vssd1
+ vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12925__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08122_ _04497_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] _04468_ team_01_WB.instance_to_wrap.cpu.f0.num\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08812__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08704__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13149__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08053_ _04512_ _04527_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08423__B net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap730 _04717_ vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_2
XFILLER_0_128_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09368__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09222__D1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15537__A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12660__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1021_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10383__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1119_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09535__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[6\] net669 _05278_ _05280_
+ _05286_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14113__A2 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout481_A _07949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08886_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[2\] net912 vssd1
+ vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__and3_1
XANTENNA__10135__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1390_A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12896__A _04837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout746_A _04682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18057__1557 vssd1 vssd1 vccd1 vccd1 _18057__1557/HI net1557 sky130_fd_sc_hd__conb_1
XANTENNA__09828__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10438__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09507_ net1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[29\] net968
+ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout913_A net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09701__C net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09438_ _05764_ _05765_ _05776_ _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09369_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[26\] _04766_ net686
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[26\] _05708_ vssd1 vssd1 vccd1
+ vccd1 _05709_ sky130_fd_sc_hd__a221o_1
XANTENNA__12835__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11400_ _04469_ _07723_ _07721_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12380_ net2219 net285 net426 vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_70 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16970__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11331_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] net1162 _04552_ _07652_ vssd1
+ vssd1 vccd1 vccd1 _07664_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17986__1486 vssd1 vssd1 vccd1 vccd1 _17986__1486/HI net1486 sky130_fd_sc_hd__conb_1
XFILLER_0_50_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08333__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14054__C _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14050_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[43\] _04256_ _04262_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[51\]
+ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__a22o_1
XANTENNA__09359__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11262_ _06135_ _06163_ _07175_ net563 vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_63_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13001_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[85\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[93\]
+ net857 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__mux2_1
X_10213_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[8\] net795 net774 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__a22o_1
XANTENNA__16200__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12570__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ _07532_ net562 _07112_ vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__and3b_1
XFILLER_0_105_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input42_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14104__A2 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[11\] net821 net778 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17740_ clknet_leaf_66_wb_clk_i _03416_ _01680_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10126__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14952_ net1276 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__inv_2
X_10075_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[7\] net971 vssd1
+ vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16350__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13903_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\] _04141_ vssd1 vssd1 vccd1 vccd1
+ _04204_ sky130_fd_sc_hd__and4_1
X_17671_ clknet_leaf_117_wb_clk_i _03356_ _01612_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14883_ net1188 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
XANTENNA__11914__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16622_ clknet_leaf_8_wb_clk_i _02309_ _00605_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13834_ net1956 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[27\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_134_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13615__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13765_ net1170 _04153_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__nand2_2
XANTENNA__13414__B _05224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16553_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[19\]
+ _00536_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10977_ net374 net342 net341 _06526_ net551 net542 vssd1 vssd1 vccd1 vccd1 _07317_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15504_ net1270 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12716_ net2851 net307 net386 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16484_ clknet_leaf_84_wb_clk_i _02238_ _00467_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13696_ _04502_ _04113_ _04117_ _04118_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__or4_2
XFILLER_0_128_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15435_ net1296 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__inv_2
X_12647_ net2606 net298 net394 vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14526__A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15366_ net1325 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__inv_2
X_12578_ net2630 net284 net401 vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08524__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17105_ clknet_leaf_15_wb_clk_i _02792_ _01088_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11529_ net1847 team_01_WB.instance_to_wrap.cpu.DM0.ihit net587 net1097 vssd1 vssd1
+ vccd1 vccd1 _03323_ sky130_fd_sc_hd__a22o_1
X_14317_ net1347 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18085_ net1585 vssd1 vssd1 vccd1 vccd1 la_data_out[127] sky130_fd_sc_hd__buf_2
X_15297_ net1249 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__inv_2
Xhold307 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18102__1589 vssd1 vssd1 vccd1 vccd1 _18102__1589/HI net1589 sky130_fd_sc_hd__conb_1
XFILLER_0_68_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10492__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold318 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
X_17036_ clknet_leaf_133_wb_clk_i _02723_ _01019_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold329 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ net1354 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__inv_2
XANTENNA__09058__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15357__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14179_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[10\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\]
+ _04448_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12480__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout809 net810 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08897__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09770__A2 _04636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17819__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ net1008 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[4\] net896 vssd1
+ vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__and3_1
Xhold1007 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[8\] vssd1 vssd1 vccd1 vccd1
+ net2623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
X_17938_ net1438 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xhold1029 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10668__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09522__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1380 net1414 vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__buf_2
Xfanout1391 net1395 vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__buf_4
X_08671_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[7\] net919 vssd1
+ vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__and3_1
X_17869_ clknet_leaf_82_wb_clk_i _03544_ _01809_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13606__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09090__A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08418__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09223_ _05554_ _05555_ _05556_ _05562_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__or4_1
XFILLER_0_107_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10840__A1 _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12655__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17923__1611 vssd1 vssd1 vccd1 vccd1 net1611 _17923__1611/LO sky130_fd_sc_hd__conb_1
XFILLER_0_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1069_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09154_ _04947_ _05492_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11396__A2 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08105_ team_01_WB.instance_to_wrap.cpu.f0.state\[2\] team_01_WB.instance_to_wrap.cpu.f0.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16223__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09085_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[13\] net883
+ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1236_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08036_ net1727 net567 net346 team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1
+ vccd1 vccd1 _03555_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold830 _02117_ vssd1 vssd1 vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 _03438_ vssd1 vssd1 vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold863 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold874 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[19\] vssd1 vssd1 vccd1 vccd1
+ net2501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1403_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold896 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[62\] vssd1 vssd1 vccd1 vccd1
+ net2512 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17499__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09987_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[2\] net803 net759 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout863_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08938_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[6\] net917 vssd1
+ vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__and3_1
Xhold1530 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3146 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10659__A1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1541 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3157 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09513__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1552 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[79\] vssd1 vssd1 vccd1 vccd1
+ net3168 sky130_fd_sc_hd__dlygate4sd3_1
X_08869_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[3\] net658 _05191_ _05192_
+ _05201_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__a2111o_1
Xhold1563 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1574 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3190 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08721__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1585 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3201 sky130_fd_sc_hd__dlygate4sd3_1
X_10900_ net517 _06969_ _07236_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__a21oi_1
X_11880_ net2662 net229 net484 vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__mux2_1
Xhold1596 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3212 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10831_ net562 _07089_ _07155_ _07170_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__a31o_2
XFILLER_0_67_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13550_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _05616_ _03925_ vssd1
+ vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__a21oi_1
X_10762_ _06945_ _07100_ net329 _06894_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12501_ net2985 net273 net409 vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10831__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13481_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _05679_ _03941_ vssd1
+ vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__a21oi_1
X_10693_ _06889_ _06907_ net538 vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__mux2_1
XANTENNA__12565__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15220_ net1267 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__inv_2
X_12432_ net3143 net206 net415 vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08344__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15151_ net1216 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__inv_2
X_12363_ net3121 net247 net424 vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14102_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[93\] _04241_ _04262_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[53\]
+ _04388_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11314_ team_01_WB.instance_to_wrap.cpu.f0.state\[3\] net1162 vssd1 vssd1 vccd1 vccd1
+ _07651_ sky130_fd_sc_hd__or2_1
X_15082_ net1272 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12294_ net2123 net221 net433 vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14033_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[82\] _04245_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[114\]
+ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__a22o_1
XANTENNA__11909__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11245_ net523 _07248_ _07584_ vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09752__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ net526 _07158_ vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__or2_1
XANTENNA__13409__B _05220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09606__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08510__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16866__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ _05301_ _06466_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__xor2_1
X_15984_ net1336 vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17723_ clknet_leaf_109_wb_clk_i _00016_ _01664_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10058_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] net627 _06396_ _06397_
+ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__a22o_2
X_14935_ net1199 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17654_ clknet_leaf_90_wb_clk_i _03339_ _01595_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14866_ net1232 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08519__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09114__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16605_ clknet_leaf_48_wb_clk_i _02292_ _00588_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13817_ net2152 net834 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[10\]
+ sky130_fd_sc_hd__and2_1
X_17585_ clknet_leaf_79_wb_clk_i _03272_ _01544_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09268__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14797_ net1212 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_69_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_85_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16536_ clknet_leaf_110_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[2\]
+ _00519_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13748_ team_01_WB.instance_to_wrap.cpu.c0.count\[3\] team_01_WB.instance_to_wrap.cpu.c0.count\[2\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[1\] vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10822__A1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12475__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16467_ clknet_leaf_141_wb_clk_i _02221_ _00450_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08491__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13679_ team_01_WB.instance_to_wrap.cpu.c0.count\[4\] team_01_WB.instance_to_wrap.cpu.c0.count\[5\]
+ _04101_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__and3_1
XANTENNA__14256__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15418_ net1192 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__inv_2
X_16398_ clknet_leaf_69_wb_clk_i _02152_ _00381_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15349_ net1219 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__inv_2
XANTENNA__09440__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold104 _02026_ vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold115 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[29\] vssd1 vssd1 vccd1 vccd1
+ net1731 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09991__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18068_ net1568 vssd1 vssd1 vccd1 vccd1 la_data_out[110] sky130_fd_sc_hd__buf_2
Xhold126 net99 vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18056__1556 vssd1 vssd1 vccd1 vccd1 _18056__1556/HI net1556 sky130_fd_sc_hd__conb_1
Xhold137 team_01_WB.instance_to_wrap.a1.ADR_I\[1\] vssd1 vssd1 vccd1 vccd1 net1753
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17641__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11819__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold148 team_01_WB.instance_to_wrap.cpu.f0.write_data\[21\] vssd1 vssd1 vccd1 vccd1
+ net1764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 net119 vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] net627 _06248_ _06249_
+ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__a22o_2
X_17019_ clknet_leaf_50_wb_clk_i _02706_ _01002_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout606 net609 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09085__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09841_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[13\] net819 net772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__a22o_1
XANTENNA__09743__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout628 _03739_ vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout639 net642 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09772_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[15\] net822 net780 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__a22o_1
XANTENNA__17791__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08723_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[5\] net914 vssd1
+ vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_52_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout277_A _07851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08654_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[10\] net879
+ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_1_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17985__1485 vssd1 vssd1 vccd1 vccd1 _17985__1485/HI net1485 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_1_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17021__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08585_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[15\] net887
+ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout444_A _07959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1186_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12385__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17171__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout611_A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1353_A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09206_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[17\] net878
+ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__and3_1
XANTENNA__16739__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09137_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[14\] net902
+ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09982__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[12\] _04776_ _05382_
+ _05400_ _05401_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_113_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout980_A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08019_ _04512_ _04514_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__nor2_1
XANTENNA__16889__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold671 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11030_ _05455_ net374 vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold682 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 _01986_ vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08330__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16119__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12981_ net1745 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[113\] net866 vssd1 vssd1
+ vccd1 vccd1 _02144_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1360 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2976 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1371 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[89\] vssd1 vssd1 vccd1 vccd1
+ net2987 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ net1316 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1382 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2998 sky130_fd_sc_hd__dlygate4sd3_1
X_11932_ net2104 net209 net477 vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__mux2_1
Xhold1393 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net3009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11863_ net2236 net218 net483 vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__mux2_1
X_14651_ net1251 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__inv_2
XANTENNA__09161__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16269__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17514__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13602_ net724 _07553_ net1067 vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__o21a_1
X_10814_ net344 _07091_ _07136_ _07153_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_67_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17370_ clknet_leaf_45_wb_clk_i _03057_ _01353_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14582_ net1390 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11794_ net2252 net221 net491 vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16321_ clknet_leaf_64_wb_clk_i _02075_ _00304_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[44\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_81_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10745_ _06906_ _07084_ net339 vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__o21a_1
X_13533_ net197 net193 _07850_ net643 vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__o211a_1
XANTENNA__12295__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13464_ _03923_ _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10280__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16252_ clknet_leaf_80_wb_clk_i net1726 _00240_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
X_10676_ _07004_ _07015_ net528 vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15203_ net1186 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__inv_2
X_12415_ net2272 net281 net420 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16183_ clknet_leaf_113_wb_clk_i _01943_ _00171_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13395_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] _04847_ vssd1 vssd1
+ vccd1 vccd1 _03856_ sky130_fd_sc_hd__xor2_1
XANTENNA__10568__A0 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12346_ net2243 net254 net427 vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15134_ net1275 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09973__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_116_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15065_ net1258 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12277_ net2555 net256 net435 vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14016_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[65\] _04233_ _04245_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[81\]
+ _04306_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11228_ _06748_ _06749_ _05967_ vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__a21o_1
XANTENNA__11532__A2 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15635__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11159_ _06928_ _07497_ _07498_ _06920_ vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__a22o_1
XANTENNA__17044__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17922__1610 vssd1 vssd1 vccd1 vccd1 net1610 _17922__1610/LO sky130_fd_sc_hd__conb_1
XANTENNA__09633__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15967_ net1409 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__inv_2
XANTENNA__10779__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17706_ clknet_leaf_101_wb_clk_i _03390_ _01647_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14918_ net1299 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15898_ net1383 vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17637_ clknet_leaf_117_wb_clk_i _03322_ _01578_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14849_ net1239 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__inv_2
X_08370_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\]
+ _04709_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__nand3_2
X_17568_ clknet_leaf_61_wb_clk_i _03255_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12796__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13993__B1 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16519_ clknet_leaf_115_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[17\]
+ _00502_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10718__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17499_ clknet_leaf_50_wb_clk_i _03186_ _01482_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10023__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__A1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09964__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11220__B2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08712__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08431__B net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09716__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout403 _03565_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_6
Xfanout414 _03563_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_4
Xfanout425 _07966_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_54_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13764__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout394_A _03568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 _07963_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09824_ _06159_ _06161_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__xnor2_2
Xfanout447 _07958_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_8
Xfanout458 _07956_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1101_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout469 net470 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_35_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_14__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09755_ _06073_ _06083_ _06084_ _06094_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13276__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout561_A _04749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[5\] net903 vssd1
+ vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08409__A_N _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09686_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[22\] net790 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[22\]
+ _06003_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08637_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[10\] net881 vssd1
+ vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08568_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[19\] net691 _04905_ _04906_
+ _04907_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_77_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16561__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17687__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12787__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13984__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08499_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ _04622_ _04719_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__nand4_2
XANTENNA__10798__A0 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10628__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10530_ _06865_ _06867_ _06869_ vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_98_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11032__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10461_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[26\] net808 _06787_
+ _06791_ _06794_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12843__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13200__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12200_ net2826 net202 net443 vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11211__A1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13180_ team_01_WB.instance_to_wrap.a1.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1
+ _03736_ sky130_fd_sc_hd__and2_1
X_10392_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[16\] net805 net744 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12131_ net2892 net209 net452 vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17067__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ net2274 net216 net459 vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__mux2_1
Xhold490 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09156__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11013_ _07142_ _07143_ _07095_ vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_70_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16870_ clknet_leaf_42_wb_clk_i _02557_ _00853_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout970 _04638_ vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__buf_2
X_15821_ net1317 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__inv_2
Xfanout981 _04499_ vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout992 net993 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_126_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15752_ net1400 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12964_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[0\] _05150_ net1036 vssd1
+ vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1190 team_01_WB.instance_to_wrap.cpu.K0.code\[7\] vssd1 vssd1 vccd1 vccd1 net2806
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08143__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16904__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14703_ net1319 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__inv_2
X_11915_ net2791 net285 net482 vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ net1186 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ net357 _03670_ _03671_ net870 net1886 vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__a32o_1
XANTENNA__08694__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11922__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18055__1555 vssd1 vssd1 vccd1 vccd1 _18055__1555/HI net1555 sky130_fd_sc_hd__conb_1
XFILLER_0_135_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17422_ clknet_leaf_8_wb_clk_i _03109_ _01405_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ net1212 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__inv_2
X_11846_ net1979 net287 net489 vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12778__A1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12778__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17353_ clknet_leaf_23_wb_clk_i _03040_ _01336_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11777_ net2313 net256 net496 vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__mux2_1
X_14565_ net1406 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16304_ clknet_leaf_73_wb_clk_i net2502 _00287_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10728_ net515 _07067_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__nand2_1
X_13516_ net197 net193 _07837_ net643 vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__o211a_1
X_17284_ clknet_leaf_51_wb_clk_i _02971_ _01267_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14496_ net1337 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16235_ clknet_leaf_105_wb_clk_i net1908 _00223_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10659_ _06158_ net374 net544 vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13447_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _05380_ vssd1 vssd1
+ vccd1 vccd1 _03908_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14534__A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10005__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ _05834_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 _03839_ sky130_fd_sc_hd__and2b_1
X_16166_ clknet_leaf_97_wb_clk_i _01929_ _00154_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17984__1484 vssd1 vssd1 vccd1 vccd1 _17984__1484/HI net1484 sky130_fd_sc_hd__conb_1
XANTENNA__12950__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15117_ net1213 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__inv_2
X_12329_ net3052 _07838_ net429 vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__mux2_1
X_16097_ clknet_leaf_83_wb_clk_i _01872_ _00085_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15048_ net1290 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__inv_2
XANTENNA__16434__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16999_ clknet_leaf_16_wb_clk_i _02686_ _00982_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_84_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_30_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09540_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[28\] _04665_
+ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09331__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09471_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[30\] net915 vssd1
+ vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11832__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08422_ net1107 net1110 net1113 net1115 vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_138_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10956__B _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08707__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08353_ _04690_ _04691_ _04692_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__or3_1
XANTENNA__12769__B2 _03607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08426__B net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10244__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11441__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08284_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__and4b_1
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12663__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1051_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout407_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09398__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1149_A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14143__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout200 _07633_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout776_A _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1209 net1210 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13497__A2 _06961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout211 net212 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_2
XFILLER_0_100_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout222 _07831_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__buf_2
XFILLER_0_100_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout233 net234 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_2
Xfanout244 _07862_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_1
XFILLER_0_22_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout255 net258 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__buf_2
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout266 _07880_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09807_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[14\] net812 net781 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__a22o_1
Xfanout277 _07851_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_2
Xfanout288 net290 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_2
Xfanout299 net301 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__buf_2
XANTENNA__09704__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout943_A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07999_ team_01_WB.instance_to_wrap.cpu.f0.num\[3\] vssd1 vssd1 vccd1 vccd1 _04497_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11308__A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[20\] net963
+ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09322__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11027__B _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12838__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[22\] net945
+ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__and3_1
XANTENNA__11742__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11700_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[11\] net717 vssd1 vssd1 vccd1
+ vccd1 _07897_ sky130_fd_sc_hd__or2_1
X_12680_ net1997 net299 net388 vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11631_ net2860 net248 net500 vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08336__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10235__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11562_ net3199 _07786_ net35 vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__a21o_1
X_14350_ net1363 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__inv_2
XANTENNA__11432__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16307__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ _06849_ _06850_ _06851_ _06852_ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__or4_1
X_13301_ net565 _03784_ net829 vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14281_ net1374 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__inv_2
XANTENNA__12573__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11493_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[16\] net579 vssd1 vssd1 vccd1
+ vccd1 _07774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13232_ net3075 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1
+ vccd1 vccd1 _01918_ sky130_fd_sc_hd__a22o_1
X_16020_ net1377 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__inv_2
XANTENNA__09928__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[26\] net972
+ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__and3_1
XANTENNA_input72_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11196__A0 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10538__A3 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13163_ net1899 net850 net841 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[13\] vssd1
+ vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10375_ _06712_ _06714_ vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__nand2_1
XANTENNA__10943__A0 _07156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08600__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17702__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08071__B _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12114_ net2694 net283 net458 vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__mux2_1
XANTENNA__14134__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17971_ net1471 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
X_13094_ _03717_ net2410 net860 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11917__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16922_ clknet_leaf_45_wb_clk_i _02609_ _00905_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12045_ net2052 net287 net465 vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__mux2_1
XANTENNA__15185__A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09183__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13417__B _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16853_ clknet_leaf_123_wb_clk_i _02540_ _00836_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17852__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15804_ net1323 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16784_ clknet_leaf_15_wb_clk_i _02471_ _00767_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13996_ _04273_ _04275_ _04277_ _04287_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__or4_2
XFILLER_0_1_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09911__A _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15735_ net1198 vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12947_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[8\] net1035 vssd1 vssd1 vccd1
+ vccd1 _03708_ sky130_fd_sc_hd__or2_1
XANTENNA__11120__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14529__A net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13660__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11671__A1 _07232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15666_ net1233 vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12878_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[29\] _03659_ net1031 vssd1
+ vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__mux2_1
XANTENNA__08527__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17405_ clknet_leaf_21_wb_clk_i _03092_ _01388_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14617_ net1360 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__inv_2
X_11829_ net2059 net220 net488 vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__mux2_1
X_15597_ net1211 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17336_ clknet_leaf_30_wb_clk_i _03023_ _01319_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11423__A1 _07701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14548_ net1392 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10777__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12483__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_131_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17267_ clknet_leaf_129_wb_clk_i _02954_ _01250_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14479_ net1332 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14264__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16218_ clknet_leaf_78_wb_clk_i net1741 _00206_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09919__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17198_ clknet_leaf_6_wb_clk_i _02885_ _01181_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16149_ clknet_leaf_96_wb_clk_i net2920 _00137_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[8\] net694 _05308_ _05309_
+ _05310_ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__a2111o_1
XANTENNA_clkbuf_leaf_109_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17725__D net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11827__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15095__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold19 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[11\] vssd1 vssd1 vccd1 vccd1
+ net1635 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09093__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09523_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[29\] net808 net748 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08658__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12658__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout357_A net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1099_A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[29\] net684 _04797_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[29\] vssd1 vssd1 vccd1 vccd1
+ _05794_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11662__A1 _07135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08405_ _04732_ _04739_ _04740_ _04742_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__and4_1
XFILLER_0_93_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09385_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[26\] net647 _05720_
+ _05721_ _05724_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_30_1502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout524_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1266_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10217__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ net1131 net948 vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_95_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08267_ net2562 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[6\] net1037 vssd1 vssd1
+ vccd1 vccd1 _03420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12393__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17725__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08198_ net2815 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[75\] net1051 vssd1 vssd1
+ vccd1 vccd1 _03489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout893_A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08043__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08594__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14116__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10160_ net341 _06497_ _06498_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__and3_1
X_18054__1554 vssd1 vssd1 vccd1 vccd1 _18054__1554/HI net1554 sky130_fd_sc_hd__conb_1
XFILLER_0_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 net1009 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1017 net1024 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__buf_2
X_10091_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[7\] net818 net807 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__a22o_1
Xfanout1028 net1029 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__buf_2
Xfanout1039 net1045 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17105__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13850_ net1166 net1060 net1798 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[11\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13627__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12801_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[9\] _07269_ net1028 vssd1 vssd1
+ vccd1 vccd1 _03629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13781_ net1170 _04160_ _04163_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__and3_1
X_10993_ _05115_ _07324_ _07332_ _07069_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_96_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10877__A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12568__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13642__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17983__1483 vssd1 vssd1 vccd1 vccd1 _17983__1483/HI net1483 sky130_fd_sc_hd__conb_1
X_15520_ net1244 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__inv_2
X_12732_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] net1054 net363 _03581_
+ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__a22o_1
XANTENNA__11653__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10456__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08347__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17255__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15451_ net1197 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12663_ net2455 net205 net387 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__mux2_1
X_14402_ net1333 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10208__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11405__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11614_ net721 _07056_ _07828_ vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__o21ai_1
X_15382_ net1223 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12594_ net2179 net248 net397 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17121_ clknet_leaf_44_wb_clk_i _02808_ _01104_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14333_ net1370 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11545_ net1623 net1158 net589 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1
+ vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17052_ clknet_leaf_32_wb_clk_i _02739_ _01035_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11476_ net368 _07765_ net2886 net874 vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__o2bb2a_1
X_14264_ net1323 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16003_ net1399 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12905__A1 _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08513__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08034__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13215_ net2 net836 net629 net3076 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__o22a_1
X_10427_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[27\] net818 net758 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14195_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[16\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\]
+ _04458_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__and3_1
X_13146_ net1703 net844 net839 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[30\] vssd1
+ vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a22o_1
X_10358_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[17\] net779 net750 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__a22o_1
XANTENNA__11647__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13077_ net2727 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[17\] net866 vssd1 vssd1
+ vccd1 vccd1 _02048_ sky130_fd_sc_hd__mux2_1
XANTENNA__10551__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17954_ net1454 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
X_10289_ net1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[19\] net951
+ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12028_ net2247 net222 net465 vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__mux2_1
X_16905_ clknet_leaf_9_wb_clk_i _02592_ _00888_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_17885_ clknet_leaf_104_wb_clk_i _03560_ _01825_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09344__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16836_ clknet_leaf_53_wb_clk_i _02523_ _00819_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12478__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16767_ clknet_leaf_7_wb_clk_i _02454_ _00750_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13979_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[32\] _04221_ _04246_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[40\]
+ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15718_ net1325 vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11644__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16698_ clknet_leaf_60_wb_clk_i _02385_ _00681_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15649_ net1249 vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__inv_2
XANTENNA__16622__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09170_ _05499_ _05503_ _05505_ _05509_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09065__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08121_ _04469_ team_01_WB.instance_to_wrap.cpu.f0.num\[26\] team_01_WB.instance_to_wrap.cpu.f0.num\[18\]
+ _04476_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__o22a_1
X_17319_ clknet_leaf_123_wb_clk_i _03006_ _01302_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10726__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08812__A2 _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08052_ _04528_ _04529_ _04527_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10027__A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09773__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08954_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[6\] net684 _05283_ _05285_
+ _05288_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1014_A _04490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08885_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[2\] net880 vssd1
+ vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout474_A _07952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13085__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12388__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout641_A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09506_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[29\] net969
+ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12832__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09437_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[28\] net681 net673 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[28\]
+ _05761_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout906_A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09368_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[26\] net681 net661 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08319_ net1131 net951 vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__and2_4
X_09299_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[22\] net934 vssd1
+ vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__and3_1
XANTENNA_60 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11330_ _07663_ net3006 _07655_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14054__D _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11261_ _06163_ _07175_ _06135_ vssd1 vssd1 vccd1 vccd1 _07601_ sky130_fd_sc_hd__o21a_1
XANTENNA__12851__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10212_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[8\] net817 net810 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[8\]
+ _06551_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__a221o_1
X_13000_ net2733 net2718 net852 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__mux2_1
XANTENNA__13560__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ _06598_ _06604_ _06742_ vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__and3_1
XANTENNA__08630__A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10143_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[11\] net812 net750 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09516__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14951_ net1325 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__inv_2
XANTENNA_input35_A gpio_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[7\] net978 vssd1
+ vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__and3_1
XANTENNA__09164__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13902_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ _04141_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\] vssd1 vssd1 vccd1 vccd1
+ _04203_ sky130_fd_sc_hd__a31o_1
X_17670_ clknet_leaf_117_wb_clk_i _03355_ _01611_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14882_ net1266 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
XANTENNA__10103__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16621_ clknet_leaf_138_wb_clk_i _02308_ _00604_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13833_ net2233 net832 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[26\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__12298__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13615__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16645__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10429__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16552_ clknet_leaf_115_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[18\]
+ _00535_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13764_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\]
+ net604 vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10400__A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10976_ _07015_ net329 _07312_ _07315_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__a22o_1
X_15503_ net1216 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__inv_2
X_12715_ net2087 net312 net384 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08508__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16483_ clknet_leaf_94_wb_clk_i _02237_ _00466_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13695_ team_01_WB.instance_to_wrap.cpu.c0.count\[11\] team_01_WB.instance_to_wrap.cpu.c0.count\[8\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[15\] team_01_WB.instance_to_wrap.cpu.c0.count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__or4bb_1
XANTENNA__11930__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15434_ net1279 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12646_ net2050 net280 net392 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16795__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08805__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12051__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15365_ net1208 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12577_ net2098 net251 net400 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17104_ clknet_leaf_128_wb_clk_i _02791_ _01087_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14316_ net1346 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__inv_2
X_11528_ net1659 net1157 net590 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1
+ vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__a22o_1
X_18084_ net1584 vssd1 vssd1 vccd1 vccd1 la_data_out[126] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15296_ net1244 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold308 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[5\] vssd1 vssd1 vccd1 vccd1
+ net1935 sky130_fd_sc_hd__dlygate4sd3_1
X_17035_ clknet_leaf_0_wb_clk_i _02722_ _01018_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14247_ net1354 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__inv_2
XANTENNA__14542__A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11459_ _04753_ _07630_ vssd1 vssd1 vccd1 vccd1 _07755_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09636__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14178_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\] _04448_ net1778 vssd1
+ vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13129_ net1725 net850 net633 team_01_WB.instance_to_wrap.a1.ADR_I\[14\] vssd1 vssd1
+ vccd1 vccd1 _02012_ sky130_fd_sc_hd__a22o_1
XANTENNA__16175__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13303__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1008 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[74\] vssd1 vssd1 vccd1 vccd1
+ net2624 sky130_fd_sc_hd__dlygate4sd3_1
X_17937_ net1437 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
Xhold1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout1370 net1379 vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__buf_4
XFILLER_0_108_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08670_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[7\] net926 vssd1
+ vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__and3_1
XANTENNA__10668__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1381 net1389 vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17868_ clknet_leaf_94_wb_clk_i _03543_ _01808_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1392 net1395 vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__buf_4
X_16819_ clknet_leaf_137_wb_clk_i _02506_ _00802_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_17799_ clknet_leaf_63_wb_clk_i _03475_ _01739_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[69\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__13606__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17570__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12001__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18053__1553 vssd1 vssd1 vccd1 vccd1 _18053__1553/HI net1553 sky130_fd_sc_hd__conb_1
XANTENNA__11840__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09222_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[17\] net691 _05544_ _05545_
+ net706 vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10840__A2 _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14031__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08715__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09153_ _04947_ _05492_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout222_A _07831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08104_ team_01_WB.instance_to_wrap.cpu.f0.state\[2\] _04563_ _04574_ vssd1 vssd1
+ vccd1 vccd1 _04575_ sky130_fd_sc_hd__and3_1
XANTENNA__10053__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09994__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09084_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[13\] net902
+ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13767__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08035_ net1789 net567 net346 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1
+ vccd1 vccd1 _03556_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold820 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12671__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1131_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold831 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1229_A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold842 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13542__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16518__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold853 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] vssd1 vssd1 vccd1 vccd1
+ net2469 sky130_fd_sc_hd__dlygate4sd3_1
X_17982__1482 vssd1 vssd1 vccd1 vccd1 _17982__1482/HI net1482 sky130_fd_sc_hd__conb_1
Xhold864 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08450__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold875 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[0\] vssd1 vssd1 vccd1 vccd1
+ net2491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 _02058_ vssd1 vssd1 vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_A _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold897 _03476_ vssd1 vssd1 vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09986_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[2\] _04684_ net771 vssd1
+ vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__a21o_1
X_08937_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[6\] net937 vssd1
+ vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout856_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11305__B1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16668__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1520 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 team_01_WB.instance_to_wrap.cpu.f0.num\[31\] vssd1 vssd1 vccd1 vccd1 net3147
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1553 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3169 sky130_fd_sc_hd__dlygate4sd3_1
X_08868_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[3\] net700 net680 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__a22o_1
Xhold1564 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1575 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[14\] vssd1 vssd1 vccd1 vccd1 net3191
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1586 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1597 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 net3213
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08799_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[0\] net935 vssd1
+ vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_64_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10830_ _07169_ _07163_ _07162_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__or3b_1
XANTENNA__11608__A1 _07019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12805__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08328__C net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10761_ net532 _06904_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__nor2_1
XANTENNA__12846__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11750__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ net2194 net243 net407 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09029__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10692_ net536 _06896_ _07031_ net376 vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__o211a_1
X_13480_ _03934_ _03936_ _03938_ _03940_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__o31a_1
XFILLER_0_137_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14022__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12431_ net3193 net274 net416 vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08344__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09985__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15150_ net1283 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12362_ net3215 net214 net424 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14101_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[69\] _04247_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[61\]
+ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15458__A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11313_ _04504_ team_01_WB.instance_to_wrap.cpu.f0.state\[3\] net585 vssd1 vssd1
+ vccd1 vccd1 _00019_ sky130_fd_sc_hd__a21o_1
XANTENNA__12581__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15081_ net1228 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__inv_2
X_12293_ net3246 net224 net431 vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16198__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13533__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14032_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[42\] _04246_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[122\]
+ _04312_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__a221o_1
X_11244_ _06906_ _06987_ _06991_ _05263_ net339 vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ net376 _06922_ _07068_ net529 vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_43_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08960__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ _05264_ _05265_ net378 vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15983_ net1405 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10418__A_N net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17722_ clknet_leaf_108_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_write_i
+ _01663_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.WRITE_I sky130_fd_sc_hd__dfrtp_2
XANTENNA__17593__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] net766 net623 vssd1
+ vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__o21a_1
X_14934_ net1201 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_82_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09191__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17653_ clknet_leaf_92_wb_clk_i _03338_ _01594_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14865_ net1292 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16604_ clknet_leaf_39_wb_clk_i _02291_ _00587_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13816_ net1672 net834 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[9\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_114_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10130__A _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17584_ clknet_leaf_80_wb_clk_i _03271_ _01543_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14796_ net1181 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16535_ clknet_leaf_108_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[1\]
+ _00518_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_70_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13747_ _04504_ team_01_WB.instance_to_wrap.cpu.DM0.state\[2\] _07783_ net3061 vssd1
+ vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__a22o_1
X_10959_ _06958_ _07101_ _07295_ _07298_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__14537__A net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10283__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16466_ clknet_leaf_122_wb_clk_i _02220_ _00449_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13678_ team_01_WB.instance_to_wrap.cpu.c0.count\[3\] team_01_WB.instance_to_wrap.cpu.c0.count\[2\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[1\] team_01_WB.instance_to_wrap.cpu.c0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__and4_1
XANTENNA__14013__A2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15417_ net1255 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_2__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12629_ net2516 net274 net393 vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__mux2_1
X_16397_ clknet_leaf_85_wb_clk_i net1833 _00380_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_38_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15348_ net1264 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__inv_2
XANTENNA__10586__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold105 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 net1721
+ sky130_fd_sc_hd__dlygate4sd3_1
X_18067_ net1567 vssd1 vssd1 vccd1 vccd1 la_data_out[109] sky130_fd_sc_hd__buf_2
XANTENNA__12491__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15279_ net1214 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold116 net98 vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold127 _02029_ vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[13\] vssd1 vssd1 vccd1 vccd1
+ net1754 sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ clknet_leaf_60_wb_clk_i _02705_ _01001_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13524__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold149 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09366__A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11535__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09840_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[13\] net805 net775 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[13\]
+ _06179_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__a221o_1
Xfanout607 net609 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout629 _03739_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__buf_2
XANTENNA__16810__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_13__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09771_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[15\] net778 net762 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[15\]
+ _06108_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11835__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08722_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[5\] net887 vssd1
+ vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08703__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[10\] net913
+ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__and3_1
XANTENNA__16960__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09532__C net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10040__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09259__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08584_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[15\] net916 vssd1
+ vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13864__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12666__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1081_A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout437_A _07963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1179_A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13351__A team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_119_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14004__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09205_ net1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[17\] net878
+ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout604_A _04151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10026__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1346_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09136_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[14\] net936 vssd1
+ vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__and3_1
XANTENNA__09967__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11223__C1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09431__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09067_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[12\] net694 _05390_ _05392_
+ _05398_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_113_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08018_ team_01_WB.instance_to_wrap.cpu.K0.code\[0\] _04513_ team_01_WB.instance_to_wrap.cpu.K0.code\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__or3b_2
XFILLER_0_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11526__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout973_A _04633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16490__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold694 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09969_ _06305_ _06306_ _06307_ _06308_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12980_ net2725 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[114\] net868 vssd1 vssd1
+ vccd1 vccd1 _02145_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1350 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1361 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[34\] vssd1 vssd1 vccd1 vccd1
+ net2977 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11931_ net2403 net248 net477 vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__mux2_1
Xhold1372 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2988 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1383 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1394 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11046__A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14650_ net1243 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11862_ net2706 net220 net485 vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13601_ net186 _04042_ _04043_ net729 vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__a211o_1
X_10813_ _07054_ _07151_ _07152_ _07148_ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_32_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14581_ net1409 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12576__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11793_ net3083 net223 net491 vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16320_ clknet_leaf_73_wb_clk_i _02074_ _00303_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13261__A _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13532_ _03939_ _03940_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_81_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10744_ _06986_ _06989_ net537 vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16251_ clknet_leaf_95_wb_clk_i net2392 _00239_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13203__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13463_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _05616_ vssd1 vssd1
+ vccd1 vccd1 _03924_ sky130_fd_sc_hd__xor2_1
X_10675_ _07009_ _07014_ net520 vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__mux2_2
XFILLER_0_84_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15202_ net1266 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12414_ net2208 net304 net420 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16182_ clknet_leaf_112_wb_clk_i _01942_ _00170_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13394_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] _04885_ vssd1 vssd1
+ vccd1 vccd1 _03855_ sky130_fd_sc_hd__and2_1
XANTENNA__10568__A1 _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09422__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15133_ net1253 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12345_ net2762 net230 net428 vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13506__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15064_ net1176 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__inv_2
X_12276_ net3042 net260 net437 vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08090__A team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14015_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[65\] _04247_ _04265_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08521__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11227_ _06748_ _06749_ _05967_ vssd1 vssd1 vccd1 vccd1 _07567_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18052__1552 vssd1 vssd1 vccd1 vccd1 _18052__1552/HI net1552 sky130_fd_sc_hd__conb_1
XFILLER_0_43_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09914__A _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11158_ net528 _07049_ _07496_ vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__a21oi_1
XANTENNA__16983__CLK clknet_leaf_137_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10109_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[6\] net804 _04678_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__a22o_1
X_15966_ net1393 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__inv_2
X_11089_ _07352_ _07422_ _07425_ _07341_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09489__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14917_ net1208 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
X_17705_ clknet_leaf_103_wb_clk_i _03389_ _01646_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_15897_ net1337 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__inv_2
XANTENNA__17339__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10498__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17636_ clknet_leaf_116_wb_clk_i _03321_ _01577_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14848_ net1244 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12486__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17567_ clknet_leaf_59_wb_clk_i _03254_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14779_ net1197 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17981__1481 vssd1 vssd1 vccd1 vccd1 _17981__1481/HI net1481 sky130_fd_sc_hd__conb_1
XANTENNA__14267__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16518_ clknet_leaf_115_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[16\]
+ _00501_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17498_ clknet_leaf_58_wb_clk_i _03185_ _01481_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17489__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16449_ clknet_leaf_54_wb_clk_i _02203_ _00432_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10008__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09413__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10559__A1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09096__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout404 _03565_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_4
XANTENNA__10035__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14730__A net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout415 _03562_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout426 _07966_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_54_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09823_ _06162_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__inv_2
Xfanout437 _07963_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_6
Xfanout448 _07958_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_4
Xfanout459 _07955_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout387_A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[20\] net783 net762 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__a22o_1
X_08705_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[5\] net880 vssd1
+ vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09685_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[22\] net811 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[22\]
+ _06006_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout554_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1296_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08636_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[10\] net888
+ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__and3_1
XANTENNA__10201__C net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12396__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[19\] net889 vssd1
+ vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__and3_1
XANTENNA__13433__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout819_A _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10247__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08498_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ _04622_ _04719_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__and4_2
XANTENNA__10798__A1 _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09652__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13736__A1 team_01_WB.instance_to_wrap.cpu.K0.keyvalid vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10460_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[26\] net789 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[26\]
+ _06799_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_115_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09404__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11252__C_N net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09119_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[14\] net911
+ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_111_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08612__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10391_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[16\] net795 net732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[16\]
+ _06717_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12130_ net2626 net248 net454 vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08341__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15736__A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ net2348 net220 net461 vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__mux2_1
XANTENNA__14640__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold480 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1
+ net2107 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09734__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ _07341_ _07347_ _07349_ _07351_ vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_70_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16236__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15820_ net1317 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__inv_2
XANTENNA__13256__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout971 _04635_ vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_5_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout982 net984 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout993 _04491_ vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__buf_4
XANTENNA__10599__B _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_137_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15751_ net1401 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__inv_2
X_12963_ net2358 net872 net359 _03716_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a22o_1
XANTENNA__09172__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11278__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13672__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1180 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2807 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ net1318 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11914_ net2138 net254 net481 vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15682_ net1260 vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16386__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12894_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[24\] net1030 vssd1 vssd1 vccd1
+ vccd1 _03671_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17421_ clknet_leaf_138_wb_clk_i _03108_ _01404_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17631__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14633_ net1184 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__inv_2
X_11845_ net3069 net257 net489 vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10238__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17352_ clknet_leaf_22_wb_clk_i _03039_ _01335_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14564_ net1393 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__inv_2
X_11776_ net2199 net259 net496 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16303_ clknet_leaf_65_wb_clk_i net2567 _00286_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13515_ _03945_ _03947_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__xor2_1
XANTENNA__08516__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17283_ clknet_leaf_21_wb_clk_i _02970_ _01266_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10727_ _06968_ _07066_ net540 vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__mux2_1
X_14495_ net1332 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16234_ clknet_leaf_105_wb_clk_i net1699 _00222_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_1
X_13446_ _03905_ _03906_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__and2_1
X_10658_ net342 net341 net544 vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08813__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16165_ clknet_leaf_99_wb_clk_i _01928_ _00153_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13377_ net1909 net830 _03838_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1
+ vccd1 vccd1 _01870_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10589_ net376 _06928_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15116_ net1209 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__inv_2
X_12328_ net3047 net216 net429 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__mux2_1
XANTENNA__12950__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16096_ clknet_leaf_83_wb_clk_i _01871_ _00084_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10961__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15047_ net1300 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__inv_2
X_12259_ net2946 net189 net435 vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__mux2_1
XANTENNA__14550__A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17161__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16998_ clknet_leaf_42_wb_clk_i _02685_ _00981_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09082__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15949_ net1411 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09470_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[30\] net931 vssd1
+ vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08421_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[23\] net934 vssd1
+ vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_138_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17619_ clknet_leaf_110_wb_clk_i _03304_ _01560_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_138_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10229__B1 _04678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11414__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12769__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08352_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[30\] net791 net788 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08283_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_138_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09819__A _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08723__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10972__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13194__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1044_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13775__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16259__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15556__A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1211_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout201 net202 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout212 _07847_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout223 net226 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_2
XFILLER_0_10_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout671_A _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 _07884_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_2
Xfanout245 net246 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_2
XANTENNA_fanout769_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout256 net258 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_2
X_09806_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[14\] net784 net732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__a22o_1
Xfanout267 net270 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_2
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10180__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout289 net290 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_2
X_07998_ team_01_WB.instance_to_wrap.cpu.f0.num\[6\] vssd1 vssd1 vccd1 vccd1 _04496_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09737_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[20\] net979
+ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout936_A _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10468__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09668_ net987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[22\] net951 vssd1
+ vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08619_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[11\] net697 net658 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__a22o_1
XANTENNA__13406__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[24\] net946 vssd1
+ vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__and3_1
XANTENNA__11324__A team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11630_ _07839_ _07841_ net611 vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18051__1551 vssd1 vssd1 vccd1 vccd1 _18051__1551/HI net1551 sky130_fd_sc_hd__conb_1
XANTENNA__11043__B _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12854__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11561_ net3115 net1168 net36 vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13300_ net1063 _07710_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10512_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[31\] net787 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14280_ net1375 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__inv_2
XANTENNA__17034__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11492_ net367 _07773_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[17\] net874
+ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_134_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09389__A1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13185__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13231_ net2833 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1
+ vccd1 vccd1 _01919_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10443_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[26\] net944
+ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__and3b_1
XFILLER_0_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11196__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08597__C1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13590__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ net1839 net849 net841 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[14\] vssd1
+ vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__a22o_1
XANTENNA_input65_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09167__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10374_ _06713_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12113_ net2149 net251 net455 vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15466__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17970_ net1470 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
X_13093_ _03716_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\] net857 vssd1 vssd1
+ vccd1 vccd1 _02032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17980__1480 vssd1 vssd1 vccd1 vccd1 _17980__1480/HI net1480 sky130_fd_sc_hd__conb_1
XANTENNA__09464__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12044_ net2232 net256 net463 vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__mux2_1
X_16921_ clknet_leaf_51_wb_clk_i _02608_ _00904_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16852_ clknet_leaf_12_wb_clk_i _02539_ _00835_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10171__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout790 _04654_ vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_85_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15803_ net1323 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16783_ clknet_leaf_143_wb_clk_i _02470_ _00766_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13995_ _04152_ _04283_ _04285_ _04286_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_66_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11933__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10459__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15734_ net1247 vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12946_ _05337_ _07757_ _03694_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11120__A1 _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09864__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15665_ net1292 vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__inv_2
XANTENNA__09630__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12877_ _05802_ net577 net361 vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_34_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17404_ clknet_leaf_39_wb_clk_i _03091_ _01387_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14616_ net1350 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__inv_2
X_11828_ net2795 net224 net487 vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__mux2_1
XANTENNA__14070__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15596_ net1185 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__inv_2
XANTENNA__09616__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17335_ clknet_leaf_139_wb_clk_i _03022_ _01318_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14547_ net1408 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__inv_2
X_11759_ net2997 net189 net495 vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14545__A net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09639__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17266_ clknet_leaf_129_wb_clk_i _02953_ _01249_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14478_ net1332 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16217_ clknet_leaf_105_wb_clk_i net1821 _00205_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13176__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13429_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\]
+ net595 vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__and3_1
X_17907__1599 vssd1 vssd1 vccd1 vccd1 net1599 _17907__1599/LO sky130_fd_sc_hd__conb_1
XANTENNA__16401__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17197_ clknet_leaf_140_wb_clk_i _02884_ _01180_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17527__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12923__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13581__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16148_ clknet_leaf_96_wb_clk_i _01911_ _00136_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08970_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[8\] net909 vssd1
+ vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16079_ clknet_leaf_103_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[1\]
+ _00067_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[1\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_100_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16551__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17677__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08355__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12004__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08107__A2 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11843__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[29\] net789 net780 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08718__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09855__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09453_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[29\] net689 net666 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__a22o_1
XANTENNA__09540__C _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout252_A _07904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10870__A0 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08404_ _04743_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09384_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[26\] net670 _05722_ _05723_
+ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__a211o_1
XANTENNA__14061__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08335_ net989 net971 vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__and2_2
XFILLER_0_69_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12674__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1161_A team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout517_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1259_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08266_ net3206 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\] net1047 vssd1 vssd1
+ vccd1 vccd1 _03421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13167__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08197_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[84\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[76\]
+ net1041 vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09240__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08043__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_105_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout886_A net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15286__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09284__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1007 net1009 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10090_ _06421_ _06427_ _06428_ _06429_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__or4_1
Xfanout1018 net1023 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1029 net1032 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11319__A team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10223__A _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12849__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11753__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ net3281 net640 net607 _03628_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13780_ _04164_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__inv_2
X_10992_ net531 _07286_ _07331_ net556 vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__a211o_1
XANTENNA__08503__C1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12731_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] _06961_ net1025 vssd1 vssd1
+ vccd1 vccd1 _03581_ sky130_fd_sc_hd__mux2_1
XANTENNA__11653__A2 _07621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08347__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15450_ net1189 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12662_ net2431 net277 net389 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14401_ net1339 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__inv_2
X_11613_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[29\] net716 net616 vssd1 vssd1
+ vccd1 vccd1 _07828_ sky130_fd_sc_hd__o21a_1
XANTENNA__12584__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15381_ net1220 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__inv_2
X_12593_ net3107 net214 net397 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17120_ clknet_leaf_30_wb_clk_i _02807_ _01103_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14332_ net1372 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11544_ net1638 net1158 net588 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1
+ vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17051_ clknet_leaf_20_wb_clk_i _02738_ _01034_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13158__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14263_ net1313 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__inv_2
X_11475_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[25\] net579 vssd1 vssd1 vccd1
+ vccd1 _07765_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16002_ net1390 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13214_ net13 net838 _03738_ net2066 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__a22o_1
XANTENNA__13563__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10426_ _06763_ _06764_ _06765_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__or3_1
X_14194_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\] _04458_ net1921 vssd1
+ vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11928__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ net1887 net844 net839 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[31\] vssd1
+ vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10357_ _06693_ _06694_ _06695_ _06696_ vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10392__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13076_ net2612 net2566 net858 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__mux2_1
X_17953_ net1453 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
X_10288_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[19\] net811 net794 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__a22o_1
XANTENNA__09729__B1_N net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16904_ clknet_leaf_31_wb_clk_i _02591_ _00887_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12027_ net1945 net226 net464 vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__mux2_1
XANTENNA__10133__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17884_ clknet_leaf_106_wb_clk_i _03559_ _01824_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10144__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09922__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16835_ clknet_leaf_21_wb_clk_i _02522_ _00818_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13444__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16766_ clknet_leaf_48_wb_clk_i _02453_ _00749_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13978_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[96\] _04244_ _04249_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10787__B net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12929_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[14\] net1035 vssd1 vssd1 vccd1
+ vccd1 _03696_ sky130_fd_sc_hd__or2_1
X_15717_ net1209 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__inv_2
X_16697_ clknet_leaf_47_wb_clk_i _02384_ _00680_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11644__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14043__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15648_ net1243 vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12494__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15579_ net1197 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08120_ _04471_ team_01_WB.instance_to_wrap.cpu.f0.num\[24\] _04495_ net1063 vssd1
+ vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__o2bb2a_1
X_17318_ clknet_leaf_41_wb_clk_i _03005_ _01301_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08704__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08051_ team_01_WB.instance_to_wrap.cpu.K0.code\[7\] team_01_WB.instance_to_wrap.cpu.K0.code\[6\]
+ team_01_WB.instance_to_wrap.cpu.K0.code\[5\] team_01_WB.instance_to_wrap.cpu.K0.code\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__or4b_2
X_17249_ clknet_leaf_48_wb_clk_i _02936_ _01232_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10308__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10907__A1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10027__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11838__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08576__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09816__B net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10383__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08953_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[6\] net680 _05267_ _05274_
+ _05275_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_102_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09535__C net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11139__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18050__1550 vssd1 vssd1 vccd1 vccd1 _18050__1550/HI net1550 sky130_fd_sc_hd__conb_1
X_08884_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] net730 _05111_ net1111 vssd1
+ vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_100_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10135__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1007_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12669__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout467_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09828__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[29\] net975
+ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout634_A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1376_A net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09436_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[28\] net659 _05775_
+ net707 vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14034__B1 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_111_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout801_A _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09367_ net600 _05705_ _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11602__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08318_ net1146 net1148 net1152 net1154 vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__and4_2
XFILLER_0_35_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09279__A _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_50 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[22\] net922 vssd1
+ vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__and3_1
XANTENNA_61 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ net2456 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[24\] net1046 vssd1 vssd1
+ vccd1 vccd1 _03438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11260_ net344 _07567_ _07590_ _07599_ vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__o31a_2
XFILLER_0_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10211_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[8\] net800 net744 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13560__A2 _07171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11191_ _07191_ _07521_ _07530_ vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10142_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[11\] net788 net768 vssd1
+ vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__a21o_1
X_14950_ net1325 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__inv_2
XANTENNA__13312__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[7\] net957 vssd1
+ vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13901_ net571 _04202_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__and2_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14881_ net1246 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
XANTENNA__12579__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16620_ clknet_leaf_116_wb_clk_i _02307_ _00603_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13832_ net1984 net831 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[25\]
+ sky130_fd_sc_hd__and2_1
X_16551_ clknet_leaf_115_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[17\]
+ _00534_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13763_ net604 vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09180__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10975_ _05301_ _06465_ net334 _07314_ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__a31o_1
X_15502_ net1285 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__inv_2
X_12714_ net3211 net297 net386 vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16482_ clknet_leaf_92_wb_clk_i _02236_ _00465_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__14025__B1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13694_ team_01_WB.instance_to_wrap.cpu.c0.count\[6\] _04116_ team_01_WB.instance_to_wrap.cpu.c0.count\[5\]
+ _04101_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__or4b_1
XFILLER_0_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15433_ net1228 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12645_ net2637 net304 net392 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10047__D1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15364_ net1238 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__inv_2
X_12576_ net2972 net229 net400 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__mux2_1
XANTENNA__09452__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17103_ clknet_leaf_144_wb_clk_i _02790_ _01086_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14315_ net1346 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__inv_2
XANTENNA__08524__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11527_ net1637 net1157 net590 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1
+ vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18083_ net1583 vssd1 vssd1 vccd1 vccd1 la_data_out[125] sky130_fd_sc_hd__buf_2
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15295_ net1257 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14823__A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10128__A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17034_ clknet_leaf_11_wb_clk_i _02721_ _01017_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold309 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
X_14246_ net1323 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__inv_2
X_11458_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[31\] net580 vssd1 vssd1 vccd1
+ vccd1 _07754_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08821__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10409_ _06107_ _06747_ _05999_ _06102_ _06103_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__o2111a_1
X_14177_ net2602 _04448_ _04450_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__o21a_1
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11389_ team_01_WB.instance_to_wrap.cpu.f0.i\[30\] _07696_ _07716_ vssd1 vssd1 vccd1
+ vccd1 _07718_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13128_ net81 net849 net634 net1771 vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_12__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__13303__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13059_ net2658 net2583 net864 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__mux2_1
X_17936_ net1436 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
Xhold1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout1360 net1362 vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__buf_4
Xfanout1371 net1379 vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__buf_2
Xfanout1382 net1389 vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__buf_4
X_17867_ clknet_leaf_82_wb_clk_i _03542_ _01807_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[6\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout1393 net1395 vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08730__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17715__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16818_ clknet_leaf_134_wb_clk_i _02505_ _00801_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17798_ clknet_leaf_57_wb_clk_i _03474_ _01738_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[68\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_89_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09090__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16749_ clknet_leaf_140_wb_clk_i _02436_ _00732_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14016__B1 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09691__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09221_ _05557_ _05558_ _05559_ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__or4_1
XFILLER_0_70_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10840__A3 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11422__A team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09099__A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ _05416_ _05454_ _05491_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08103_ _04568_ _04571_ _04572_ _04573_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__or4_4
XANTENNA__08434__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08797__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[13\] net933
+ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12952__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10038__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_A _07838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08034_ net1764 net568 net346 team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1
+ vccd1 vccd1 _03557_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput70 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold810 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold821 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[66\] vssd1 vssd1 vccd1 vccd1
+ net2437 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold832 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 net2459
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08549__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold854 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[50\] vssd1 vssd1 vccd1 vccd1
+ net2481 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08450__B net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1124_A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10356__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold876 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17245__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold898 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[2\] net808 net734 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08936_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[6\] net895 vssd1
+ vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__and3_1
XANTENNA__10108__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1510 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3126 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10204__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1521 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3137 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09562__A _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08867_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[3\] net927 vssd1
+ vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__and3_1
XANTENNA__12399__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1532 _01931_ vssd1 vssd1 vccd1 vccd1 net3148 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout751_A _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1543 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net3159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1554 team_01_WB.instance_to_wrap.cpu.K0.code\[1\] vssd1 vssd1 vccd1 vccd1 net3170
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout849_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1565 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08721__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1576 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3192 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10501__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08798_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[0\] net935 vssd1
+ vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__and3_1
Xhold1587 team_01_WB.instance_to_wrap.a1.ADR_I\[27\] vssd1 vssd1 vccd1 vccd1 net3203
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1598 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12805__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10816__A0 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10760_ net524 _06904_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__nor2_2
XANTENNA__14007__B1 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09682__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08906__A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09419_ _05758_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__inv_2
X_10691_ net533 _06908_ vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12430_ net2708 net211 net416 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13230__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11241__A0 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08788__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12361_ net2371 net218 net423 vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12862__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14100_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[13\] _04226_ _04259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[21\]
+ _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11312_ net830 _07649_ vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__or2_2
X_15080_ net1276 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12292_ net2939 net189 net431 vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__mux2_1
X_14031_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[66\] _04247_ _04262_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[50\]
+ _04310_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11243_ _06966_ _07527_ _06964_ vssd1 vssd1 vccd1 vccd1 _07583_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13259__A team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13533__A2 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11544__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11174_ net371 _07511_ _07513_ _06216_ _05417_ vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__o32a_1
XANTENNA__08960__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ net506 _06464_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] net627
+ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17738__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15982_ net1391 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09472__A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17721_ clknet_leaf_108_wb_clk_i _00015_ _01662_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10056_ _06384_ _06385_ _06390_ _06395_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__or4_4
X_14933_ net1220 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12102__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ clknet_leaf_92_wb_clk_i _03337_ _01593_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14864_ net1223 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__inv_2
XANTENNA__10411__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16603_ clknet_leaf_49_wb_clk_i _02290_ _00586_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08519__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13815_ net2424 net834 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[8\]
+ sky130_fd_sc_hd__and2_1
X_17583_ clknet_leaf_72_wb_clk_i _03270_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.lcd_rs
+ sky130_fd_sc_hd__dfxtp_1
X_14795_ net1295 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11941__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09268__A3 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10807__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16534_ clknet_leaf_109_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[0\]
+ _00517_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_13746_ team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] _03579_ _04137_ team_01_WB.instance_to_wrap.cpu.RU0.next_dhit
+ net834 vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__a311o_1
XFILLER_0_58_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10958_ _05042_ _06924_ _07297_ net369 vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13441__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13677_ team_01_WB.instance_to_wrap.cpu.c0.count\[1\] team_01_WB.instance_to_wrap.cpu.c0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__nand2_1
X_16465_ clknet_leaf_127_wb_clk_i _02219_ _00448_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10889_ _07017_ _07217_ _07218_ _07100_ _07226_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15416_ net1178 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__inv_2
X_12628_ net2206 net210 net393 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__mux2_1
X_16396_ clknet_leaf_77_wb_clk_i net2943 _00379_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09425__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15347_ net1278 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__inv_2
XANTENNA__15649__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12559_ net2978 net217 net401 vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14553__A net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10586__A2 _06882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16142__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15278_ net1284 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17268__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18066_ net1566 vssd1 vssd1 vccd1 vccd1 la_data_out[108] sky130_fd_sc_hd__buf_2
Xhold106 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[10\] vssd1 vssd1 vccd1 vccd1
+ net1722 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold117 _02028_ vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08551__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
X_17017_ clknet_leaf_47_wb_clk_i _02704_ _01000_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14229_ net2141 vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13524__A2 _07588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_78_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09366__B _05704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11535__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout608 net609 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__buf_2
XANTENNA__09085__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout619 _04846_ vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08951__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09770_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[15\] _04636_ net809
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[15\] vssd1 vssd1 vccd1 vccd1
+ _06110_ sky130_fd_sc_hd__a22o_1
XANTENNA__13288__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08721_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[5\] net699 net671 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__a22o_1
X_17919_ net1607 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XANTENNA__11299__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1190 net1194 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__buf_4
XANTENNA__08703__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[10\] net920
+ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__and3_1
XANTENNA__12012__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10321__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10510__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08429__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08583_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[15\] net898
+ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11851__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12799__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13460__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1074_A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09204_ net1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[17\] net931
+ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13778__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09135_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[14\] net939
+ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__and3_1
XANTENNA__12682__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1241_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1339_A net1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[12\] net671 _05389_ _05393_
+ _05397_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08461__A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout799_A _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ team_01_WB.instance_to_wrap.cpu.K0.code\[3\] team_01_WB.instance_to_wrap.cpu.K0.code\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold640 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16635__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold651 team_01_WB.instance_to_wrap.cpu.c0.count\[12\] vssd1 vssd1 vccd1 vccd1 net2267
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11526__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold673 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[50\] vssd1 vssd1 vccd1 vccd1
+ net2300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold695 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11168__A_N _07323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout966_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13807__A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09968_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[3\] net763 net751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__a22o_1
X_08919_ net602 _05224_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__nor2_1
XANTENNA__16785__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_83_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09899_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[5\] net813 _06227_ _06232_
+ _06233_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_77_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1340 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1351 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2967 sky130_fd_sc_hd__dlygate4sd3_1
X_11930_ net2745 net215 net477 vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1362 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1373 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2989 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1384 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1395 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net3011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08339__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11046__B _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ net2061 net225 net483 vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12857__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14638__A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11761__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13600_ net198 net194 _07891_ net644 vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__o211a_1
X_10812_ net555 _07141_ _07017_ vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14580_ net1393 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11792_ net2649 net190 net492 vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__mux2_1
XANTENNA__13451__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13451__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13531_ _03984_ _03985_ net1066 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\]
+ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_81_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10743_ _06990_ _06994_ net537 vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16250_ clknet_leaf_96_wb_clk_i net2034 _00238_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13462_ _03855_ _03921_ _03853_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__o21a_1
XFILLER_0_125_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10674_ _07011_ _07013_ net541 vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__mux2_2
XANTENNA__09407__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15201_ net1250 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12413_ net2792 net283 net421 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16181_ clknet_leaf_112_wb_clk_i _01941_ _00169_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13393_ _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__inv_2
XANTENNA__12592__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12962__A0 team_01_WB.instance_to_wrap.cpu.f0.write_data\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15132_ net1173 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__inv_2
X_12344_ net2344 net289 net429 vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08802__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13506__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15063_ net1200 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12275_ net3080 net233 net437 vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__mux2_1
XANTENNA__17560__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11517__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14014_ _04301_ _04302_ _04303_ _04304_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__or4_1
XANTENNA__09186__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11226_ net562 _07556_ _07557_ _07565_ vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__a31o_2
XFILLER_0_124_1680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11936__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ net527 _07025_ _07496_ vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10108_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[6\] net763 _06446_ _06447_
+ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__a211o_1
X_15965_ net1408 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__inv_2
XANTENNA__09633__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11088_ _07340_ _07427_ vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17704_ clknet_leaf_101_wb_clk_i _03388_ _01645_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_10039_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[0\] net967 vssd1
+ vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__and3_1
X_14916_ net1239 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__inv_2
XANTENNA__09894__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15896_ net1330 vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17635_ clknet_leaf_117_wb_clk_i _03320_ _01576_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_14847_ net1256 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_125_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11671__S net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17566_ clknet_leaf_61_wb_clk_i _03253_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14778_ net1192 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09110__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16517_ clknet_leaf_111_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[15\]
+ _00500_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11453__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_129_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13993__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13729_ team_01_WB.instance_to_wrap.cpu.DM0.state\[1\] team_01_WB.instance_to_wrap.cpu.DM0.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__or2_1
X_17497_ clknet_leaf_58_wb_clk_i _03184_ _01480_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_128_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16448_ clknet_leaf_19_wb_clk_i _02202_ _00431_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15379__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11205__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16379_ clknet_leaf_85_wb_clk_i _02133_ _00362_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16658__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11756__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12953__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08712__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18049_ net1549 vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__buf_2
XANTENNA__10316__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12007__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09031__D1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout405 _03565_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout416 _03562_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_4
X_09822_ _06159_ _06161_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__or2_1
XANTENNA__11846__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout427 _07965_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_54_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout438 _07963_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout449 _07958_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_8
XANTENNA__16003__A net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09753_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[20\] net733 _06090_ _06091_
+ _06092_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout282_A _07917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[5\] net911 vssd1
+ vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__and3_1
XANTENNA__09334__C1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13130__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09684_ _06020_ _06021_ _06022_ _06023_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08635_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[10\] net930 vssd1
+ vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12677__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout547_A _05152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1191_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1289_A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16188__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08566_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[19\] net886 vssd1
+ vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13433__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13984__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08497_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] net702 _04834_ _04836_
+ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__o22a_4
XFILLER_0_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11995__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13197__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09118_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[14\] _04810_
+ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10390_ _06718_ _06721_ _06726_ _06729_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__or4_1
XFILLER_0_115_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09049_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[12\] net933 vssd1
+ vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10226__A _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12060_ net2436 net225 net459 vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold470 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08376__B1 _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12172__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold492 team_01_WB.instance_to_wrap.a1.ADR_I\[30\] vssd1 vssd1 vccd1 vccd1 net2108
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11011_ _05681_ net511 vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08915__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout950 _04660_ vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__clkbuf_8
Xfanout983 net984 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13121__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout994 net996 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[1\] _05187_ net1035 vssd1
+ vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__mux2_1
XANTENNA__09876__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15750_ net1401 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__inv_2
Xhold1170 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[49\] vssd1 vssd1 vccd1 vccd1
+ net2786 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1181 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2797 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ net3129 net229 net481 vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__mux2_1
X_14701_ net1318 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__inv_2
Xhold1192 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2808 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12587__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15681_ net1240 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__inv_2
X_12893_ net362 _03669_ net1025 vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_83_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ clknet_leaf_130_wb_clk_i _03107_ _01403_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13272__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11844_ net3175 net260 net489 vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__mux2_1
X_14632_ net1296 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09628__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ net1412 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11435__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17351_ clknet_leaf_54_wb_clk_i _03038_ _01334_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11775_ net2541 net233 net497 vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11986__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08085__B _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16302_ clknet_leaf_68_wb_clk_i net2876 _00285_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13514_ net981 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] _03970_ _03971_
+ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a22o_1
X_10726_ net513 _05898_ net549 vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__mux2_1
X_17282_ clknet_leaf_36_wb_clk_i _02969_ _01265_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14494_ net1329 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13188__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16233_ clknet_leaf_104_wb_clk_i net1860 _00221_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
XANTENNA__15199__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13445_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] _05419_ vssd1 vssd1
+ vccd1 vccd1 _03906_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10657_ _06995_ _06996_ _06981_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_84_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09197__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13376_ net1834 net830 _03838_ team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1
+ vccd1 vccd1 _01871_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16164_ clknet_leaf_101_wb_clk_i _01927_ _00152_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09800__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10588_ _06900_ _06910_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__nor2_4
XANTENNA__16950__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15115_ net1297 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__inv_2
X_12327_ net2421 net222 net429 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__mux2_1
X_16095_ clknet_leaf_83_wb_clk_i _01870_ _00083_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10961__A2 _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15046_ net1290 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__inv_2
XANTENNA__09159__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12258_ _07793_ _07794_ net573 vssd1 vssd1 vccd1 vccd1 _07963_ sky130_fd_sc_hd__and3_4
XANTENNA__11666__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ net524 _07495_ vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__or2_1
XANTENNA__13854__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13447__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10174__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12189_ net2210 _07941_ net449 vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16997_ clknet_leaf_31_wb_clk_i _02684_ _00980_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13112__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09316__C1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15948_ net1387 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13663__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16330__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10477__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09660__A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09331__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12497__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15879_ net1397 vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08420_ net1006 net935 vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_138_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17618_ clknet_leaf_110_wb_clk_i _03303_ _01559_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_138_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08707__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08351_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[30\] net811 _04642_ _04644_
+ _04689_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17549_ clknet_leaf_140_wb_clk_i _03236_ _01532_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire884_A _04803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08282_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_43_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13179__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_93_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11729__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09398__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_93_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09538__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14128__C1 _04152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12960__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1037_A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14143__A2 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout497_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 net204 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_2
Xfanout213 net214 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_2
Xfanout224 net226 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10165__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout235 net238 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1204_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout246 _07862_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_2
X_09805_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[14\] net786 net769 vssd1
+ vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__a21o_1
Xfanout257 net258 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout268 net269 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_2
X_07997_ team_01_WB.instance_to_wrap.cpu.f0.num\[22\] vssd1 vssd1 vccd1 vccd1 _04495_
+ sky130_fd_sc_hd__inv_2
Xfanout279 net280 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_2
XANTENNA_fanout664_A _04806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09736_ net992 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[20\] net974 vssd1
+ vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__and3_1
XANTENNA__13654__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09322__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[22\] net975
+ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout831_A team_01_WB.instance_to_wrap.cpu.RU0.next_ihit vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08618_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[11\] net687 net648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[11\]
+ _04950_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__a221o_1
XANTENNA__16823__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11605__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12200__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[24\] net979
+ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__and3_1
XANTENNA__13406__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08549_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[19\] net694 _04886_ _04887_
+ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11324__B team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11560_ net2806 net1168 net37 vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__a21o_1
XANTENNA__11432__A3 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16973__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10511_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[31\] net772 net741 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11491_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[17\] net579 vssd1 vssd1 vccd1
+ vccd1 _07773_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13230_ net2798 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1
+ vccd1 vccd1 _01920_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09389__A2 _05726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10442_ net504 _06780_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08597__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13161_ net1723 net845 net839 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[15\] vssd1
+ vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__a22o_1
XANTENNA__16203__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13877__A_N team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10373_ _06710_ _06711_ _06708_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__o21a_1
XANTENNA__17329__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12112_ net3090 net230 net457 vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14134__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ _03715_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] net856 vssd1 vssd1
+ vccd1 vccd1 _02033_ sky130_fd_sc_hd__mux2_1
XANTENNA_input58_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12043_ net2648 net259 net463 vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__mux2_1
X_16920_ clknet_leaf_25_wb_clk_i _02607_ _00903_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09464__B _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17479__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16851_ clknet_leaf_135_wb_clk_i _02538_ _00834_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09183__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout780 net781 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__buf_6
Xfanout791 net793 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15802_ net1323 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_14__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16782_ clknet_leaf_5_wb_clk_i _02469_ _00765_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13994_ _04229_ _04238_ _04247_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[64\]
+ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09849__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ net1220 vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ net360 _03705_ _03706_ net873 net1955 vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a32o_1
XFILLER_0_133_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11120__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12110__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15664_ net1273 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12876_ net2422 net870 net357 _03658_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17403_ clknet_leaf_17_wb_clk_i _03090_ _01386_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08527__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14615_ net1360 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__inv_2
X_11827_ net3190 net189 net487 vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__mux2_1
X_15595_ net1300 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17334_ clknet_leaf_1_wb_clk_i _03021_ _01317_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14546_ net1394 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__inv_2
X_11758_ net576 _07794_ _07942_ vssd1 vssd1 vccd1 vccd1 _07943_ sky130_fd_sc_hd__and3_1
X_10709_ net515 _07024_ _06967_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_70_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17265_ clknet_leaf_15_wb_clk_i _02952_ _01248_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11689_ net2924 net260 net501 vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__mux2_1
X_14477_ net1405 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16216_ clknet_leaf_62_wb_clk_i net1853 _00204_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfrtp_1
X_13428_ _03887_ _03888_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__or2_1
X_17196_ clknet_leaf_134_wb_clk_i _02883_ _01179_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12384__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08588__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16147_ clknet_leaf_98_wb_clk_i _01910_ _00135_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13359_ net1730 _03830_ net826 vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10395__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10934__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16078_ clknet_leaf_102_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[0\]
+ _00066_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13177__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15029_ net1221 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__inv_2
XANTENNA__10147__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09552__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_140_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_140_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16846__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_1
XFILLER_0_39_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10032__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09521_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[29\] net822 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[29\]
+ _05848_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09304__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09452_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[29\] net686 net679 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[29\]
+ _05785_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__a221o_1
XANTENNA__11425__A team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12020__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08403_ _04732_ _04739_ _04742_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__nand3_2
XANTENNA__08437__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10870__A1 _06636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09383_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[26\] net699 net680 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08334_ net988 net962 vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__and2_4
XFILLER_0_35_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08265_ net2007 net2238 net1046 vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__mux2_1
XANTENNA__16226__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout412_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1154_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08196_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[85\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[77\]
+ net1039 vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12690__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08043__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14116__A2 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08594__A3 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17621__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12127__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08900__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_A _04810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1008 net1009 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_7_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1019 net1023 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09543__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11319__B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13627__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ _06055_ _06056_ _06057_ _06058_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__or4_1
X_10991_ net376 _07326_ _07328_ _07330_ _06905_ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__a32o_1
XFILLER_0_96_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09731__C net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11102__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12730_ _04510_ _03579_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__nor2_2
XFILLER_0_35_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12661_ net2217 net210 net388 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__mux2_1
XANTENNA__12865__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14400_ net1403 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11612_ net1926 net224 net499 vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12592_ net2296 net218 net397 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__mux2_1
X_15380_ net1263 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ net1688 net1158 net588 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1
+ vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14331_ net1370 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17050_ clknet_leaf_60_wb_clk_i _02737_ _01033_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14262_ net1311 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11474_ net368 _07764_ net1705 net874 vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__16719__CLK clknet_leaf_143_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16001_ net1338 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__inv_2
X_13213_ net24 net838 _03738_ net3128 vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10425_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[27\] net801 net754 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14193_ net2746 _04458_ _04460_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__o21a_1
XANTENNA__08034__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13144_ team_01_WB.instance_to_wrap.a1.curr_state\[1\] _04509_ team_01_WB.instance_to_wrap.a1.curr_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__and3b_1
XANTENNA__09475__A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10356_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[17\] net811 _06678_ _06687_
+ _06688_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09782__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_13075_ net2681 net2501 net864 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__mux2_1
X_17952_ net1452 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
XANTENNA__10414__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10287_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[19\] net807 net756 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__a22o_1
XANTENNA__12105__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12026_ net2354 net189 net464 vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__mux2_1
X_16903_ clknet_leaf_16_wb_clk_i _02590_ _00886_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_17883_ clknet_leaf_109_wb_clk_i _03558_ _01823_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11944__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16834_ clknet_leaf_34_wb_clk_i _02521_ _00817_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13618__A1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16765_ clknet_leaf_49_wb_clk_i _02452_ _00748_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13977_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[80\] _04251_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15716_ net1191 vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12928_ _05490_ _07757_ _03694_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__o21ai_1
X_16696_ clknet_leaf_27_wb_clk_i _02383_ _00679_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15647_ net1255 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__inv_2
XANTENNA__16249__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12859_ net2337 net301 net381 vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__mux2_1
XANTENNA__14043__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15578_ net1192 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__inv_2
XANTENNA__08554__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17317_ clknet_leaf_39_wb_clk_i _03004_ _01300_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14529_ net1399 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08050_ team_01_WB.instance_to_wrap.cpu.K0.code\[7\] team_01_WB.instance_to_wrap.cpu.K0.code\[5\]
+ team_01_WB.instance_to_wrap.cpu.K0.code\[4\] team_01_WB.instance_to_wrap.cpu.K0.code\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__or4b_2
XFILLER_0_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17248_ clknet_leaf_32_wb_clk_i _02935_ _01231_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09088__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17644__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap711 _04729_ vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_1
X_17179_ clknet_leaf_17_wb_clk_i _02866_ _01162_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09773__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13306__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08952_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[6\] net690 _05269_ _05276_
+ _05277_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12015__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10324__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17794__CLK clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11283__D_N _07600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11139__B _06924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08883_ _04755_ _05219_ _05221_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout195_A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11854__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13609__A1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09504_ net1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[29\] net944
+ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12832__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09435_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[28\] net697 net664 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12685__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17174__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1369_A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09366_ net598 _05704_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__or2_1
XANTENNA__08464__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08317_ net1132 net953 vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09297_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[22\] net926 vssd1
+ vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__and3_1
XANTENNA_40 _07900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_51 net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ net2587 net2353 net1050 vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout996_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15297__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08179_ net2592 net2517 net1042 vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10359__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12899__A2 _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10210_ _06547_ _06548_ _06549_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09295__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ net330 _07526_ _07529_ net556 _07525_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__a221o_1
X_10141_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[11\] net815 net779 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput180 net180 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XANTENNA__09516__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[7\] net975 vssd1
+ vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__and3_1
XANTENNA__08724__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13900_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] _04201_ vssd1 vssd1 vccd1
+ vccd1 _04202_ sky130_fd_sc_hd__xnor2_1
X_14880_ net1241 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
XANTENNA__08639__A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10531__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13831_ net2198 net831 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[24\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_97_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17517__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16550_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[16\]
+ _00533_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13762_ _04141_ _04148_ _04149_ _04150_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__and4_2
X_10974_ _05301_ net333 _07313_ net338 net371 vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15501_ net1208 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__inv_2
X_12713_ net2674 net298 net386 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__mux2_1
X_16481_ clknet_leaf_96_wb_clk_i _02235_ _00464_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12595__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13693_ team_01_WB.instance_to_wrap.cpu.c0.count\[7\] team_01_WB.instance_to_wrap.cpu.c0.count\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15432_ net1287 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12644_ net2962 net283 net393 vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__mux2_1
XANTENNA__08374__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16541__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17667__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08805__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12575_ net2573 net288 net402 vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__mux2_1
X_15363_ net1175 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17102_ clknet_leaf_6_wb_clk_i _02789_ _01085_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14314_ net1350 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11526_ net1700 team_01_WB.instance_to_wrap.cpu.DM0.ihit net587 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__a22o_1
X_18082_ net1582 vssd1 vssd1 vccd1 vccd1 la_data_out[124] sky130_fd_sc_hd__buf_2
X_15294_ net1251 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11939__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17033_ clknet_leaf_11_wb_clk_i _02720_ _01016_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10843__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ _04712_ _04753_ vssd1 vssd1 vccd1 vccd1 _07753_ sky130_fd_sc_hd__or2_1
X_14245_ net1331 vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10408_ _06598_ _06604_ _06743_ _06107_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__a211o_1
X_14176_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\] _04448_ net1412 vssd1
+ vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__a21oi_1
X_11388_ team_01_WB.instance_to_wrap.cpu.f0.i\[30\] _07716_ _07699_ vssd1 vssd1 vccd1
+ vccd1 _07717_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09636__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10339_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[17\] net958
+ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__and3_1
X_13127_ net82 net847 net632 net1712 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17047__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13058_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[28\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[36\]
+ net856 vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__mux2_1
X_17935_ team_01_WB.instance_to_wrap.cpu.LCD0.lcd_rs vssd1 vssd1 vccd1 vccd1 net157
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11674__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1350 net1351 vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__buf_4
X_12009_ net2964 net231 net469 vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__mux2_1
Xfanout1361 net1362 vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__buf_4
X_17866_ clknet_leaf_83_wb_clk_i _03541_ _01806_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_94_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1372 net1379 vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__buf_4
Xfanout1383 net1384 vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__buf_4
Xfanout1394 net1395 vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__buf_4
XFILLER_0_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16817_ clknet_leaf_19_wb_clk_i _02504_ _00800_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17797_ clknet_leaf_72_wb_clk_i _03473_ _01737_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17197__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16748_ clknet_leaf_133_wb_clk_i _02435_ _00731_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap961_A _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09691__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16679_ clknet_leaf_16_wb_clk_i _02366_ _00662_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09220_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[17\] net665 _05533_
+ _05543_ _05549_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_31_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08715__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09151_ _05456_ _05490_ net602 vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08102_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[12\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[15\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[14\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__or4b_1
XFILLER_0_126_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09082_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[13\] net935 vssd1
+ vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__and3_1
XANTENNA__10053__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09994__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11849__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08033_ net1716 net568 net346 net1063 vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold800 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
Xinput60 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold811 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
XANTENNA__16006__A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout208_A _07855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold822 _03472_ vssd1 vssd1 vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09746__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold833 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 _03456_ vssd1 vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11553__A2 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold877 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ _06318_ _06321_ _06322_ _06323_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__or4_1
Xhold899 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1117_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08935_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[6\] net890 vssd1
+ vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_73_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11305__A2 _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1500 team_01_WB.instance_to_wrap.cpu.f0.num\[13\] vssd1 vssd1 vccd1 vccd1 net3116
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1511 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3138 sky130_fd_sc_hd__dlygate4sd3_1
X_08866_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[3\] net932 vssd1
+ vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__and3_1
Xhold1533 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[55\] vssd1 vssd1 vccd1 vccd1
+ net3149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1544 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1555 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1566 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[23\] vssd1 vssd1 vccd1 vccd1
+ net3182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08797_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[0\] net691 _05134_ _05135_
+ _05136_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__a2111o_1
Xhold1577 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3193 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09281__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout744_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1588 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[87\] vssd1 vssd1 vccd1 vccd1
+ net3204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1599 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16564__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10816__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout911_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10292__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ _05756_ _05757_ net598 vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__mux2_2
X_10690_ net523 _07029_ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09349_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[25\] net681 net678 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[25\]
+ _05688_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10044__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12360_ net2013 net222 net423 vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__mux2_1
XANTENNA__11241__A1 _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09985__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08922__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11759__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11311_ _04505_ _04524_ vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12291_ _07794_ _07942_ net574 vssd1 vssd1 vccd1 vccd1 _07964_ sky130_fd_sc_hd__and3_1
X_14030_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[34\] _04230_ _04236_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[50\]
+ _04311_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_1552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11242_ _05729_ net331 _07581_ net369 vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13259__B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12741__A1 _07088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11173_ _05417_ net342 net334 _07512_ vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10124_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] net766 net623 vssd1
+ vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input40_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15981_ net1407 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17720_ clknet_leaf_109_wb_clk_i _00005_ _01661_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10055_ _06391_ _06392_ _06393_ _06394_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__or4_1
X_14932_ net1291 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
XANTENNA__10504__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09370__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ clknet_leaf_83_wb_clk_i _03336_ _01592_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14863_ net1215 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
XANTENNA__09191__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16602_ clknet_leaf_59_wb_clk_i _02289_ _00585_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13814_ net3286 net833 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[7\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_54_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17582_ clknet_leaf_77_wb_clk_i _03269_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dfxtp_1
X_14794_ net1282 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16533_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[31\]
+ _00516_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13745_ net1165 team_01_WB.instance_to_wrap.cpu.RU0.state\[2\] vssd1 vssd1 vccd1
+ vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_ihit sky130_fd_sc_hd__and2b_2
X_10957_ _06912_ _06919_ _07296_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16464_ clknet_leaf_135_wb_clk_i _02218_ _00447_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10283__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_118_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13676_ net1781 net570 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1
+ vccd1 vccd1 _01826_ sky130_fd_sc_hd__a22o_1
X_10888_ net528 _07227_ _07213_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15415_ net1201 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__inv_2
X_12627_ net2936 net249 net393 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16395_ clknet_leaf_86_wb_clk_i net2915 _00378_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15346_ net1231 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12558_ net2945 net221 net401 vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_130_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08832__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13509__B1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10586__A3 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11669__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18065_ net1565 vssd1 vssd1 vccd1 vccd1 la_data_out[107] sky130_fd_sc_hd__buf_2
X_11509_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[8\] _07756_ vssd1 vssd1 vccd1
+ vccd1 _07782_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_130_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15277_ net1207 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold107 net114 vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ _07945_ _07951_ net573 vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_130_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold118 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1
+ net1734 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold129 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[105\] vssd1 vssd1 vccd1 vccd1
+ net1745 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14182__B1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17016_ clknet_leaf_27_wb_clk_i _02703_ _00999_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_1648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14228_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] vssd1 vssd1 vccd1
+ vccd1 _02259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11535__A2 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12732__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14159_ _04187_ _04439_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout609 _03583_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09663__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08720_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[5\] net684 net680 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11299__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17918_ net1606 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_47_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09361__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1180 net1182 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__buf_4
X_08651_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[10\] net913 vssd1
+ vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__and3_1
Xfanout1191 net1194 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17849_ clknet_leaf_76_wb_clk_i net2537 _01789_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08582_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[15\] net880
+ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__and3_1
XANTENNA__10040__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12799__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09203_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[17\] net915
+ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09416__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout325_A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09134_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[14\] net928 vssd1
+ vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1067_A team_01_WB.instance_to_wrap.cpu.IM0.pc_enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09967__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11223__B2 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08742__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11579__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09065_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[12\] net667 _05388_
+ _05396_ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_60_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1234_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08461__B net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08016_ team_01_WB.instance_to_wrap.cpu.K0.code\[6\] team_01_WB.instance_to_wrap.cpu.K0.code\[5\]
+ team_01_WB.instance_to_wrap.cpu.K0.code\[4\] team_01_WB.instance_to_wrap.cpu.K0.code\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_113_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold630 _03496_ vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout694_A _04771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold641 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11526__A2 team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold663 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17362__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold674 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1401_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold696 team_01_WB.instance_to_wrap.cpu.f0.num\[1\] vssd1 vssd1 vccd1 vccd1 net2312
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09573__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09967_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[3\] net809 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout861_A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout959_A _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08918_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] net705 _05253_ _05257_
+ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__o22a_2
XANTENNA__12203__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[5\] net734 _06222_ _06226_
+ _06230_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__a2111o_1
Xhold1330 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1341 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09352__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1352 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2968 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ net599 _05187_ _05188_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__o21ai_4
Xhold1363 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2979 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1374 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1385 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[29\] vssd1 vssd1 vccd1 vccd1
+ net3001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1396 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3012 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11860_ net2933 net191 net483 vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13987__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10811_ _06969_ _07150_ _07140_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10658__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11791_ _07790_ net575 _07794_ vssd1 vssd1 vccd1 vccd1 _07944_ sky130_fd_sc_hd__and3_4
XANTENNA__09655__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11343__A team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13530_ net722 net278 net1066 vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__o21a_1
XANTENNA__11462__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10742_ _07080_ _07081_ net514 vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10673_ net550 _06340_ _07012_ vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13461_ _03854_ _03855_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nor2_1
XANTENNA__13203__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ net1237 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__inv_2
X_12412_ net2474 net253 net420 vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__mux2_1
XANTENNA__10017__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09958__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16180_ clknet_leaf_112_wb_clk_i _01940_ _00168_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13392_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] _04885_ vssd1 vssd1
+ vccd1 vccd1 _03853_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12962__A1 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15131_ net1184 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12343_ net2214 net256 net428 vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
XANTENNA__08091__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12274_ net2794 net263 net435 vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__mux2_1
X_15062_ net1202 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14013_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[41\] _04256_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[121\]
+ _04291_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__a221o_1
X_11225_ _06934_ _07201_ _07562_ _07564_ vssd1 vssd1 vccd1 vccd1 _07565_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_75_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09591__B1 _05929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11156_ net528 _07495_ vssd1 vssd1 vccd1 vccd1 _07496_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10107_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[6\] net781 net742 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__a22o_1
XANTENNA__12113__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15964_ net1387 vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__inv_2
XANTENNA__10422__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11087_ _05781_ _05899_ _07045_ _07426_ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__a31o_1
X_17703_ clknet_leaf_101_wb_clk_i _03387_ _01644_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_10038_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[0\] net953 vssd1
+ vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__and3_1
X_14915_ net1187 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15895_ net1409 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08697__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11952__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17634_ clknet_leaf_117_wb_clk_i _03319_ _01575_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14846_ net1270 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13978__B1 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17565_ clknet_leaf_59_wb_clk_i _03252_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14777_ net1306 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__inv_2
X_11989_ net2742 net319 net474 vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16516_ clknet_leaf_111_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[14\]
+ _00499_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13728_ net1156 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] team_01_WB.instance_to_wrap.cpu.DM0.enable
+ _04711_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__or4_1
XANTENNA__11453__A1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17496_ clknet_leaf_29_wb_clk_i _03183_ _01479_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16447_ clknet_leaf_35_wb_clk_i _02201_ _00430_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13659_ net727 net322 net982 vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10008__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11205__A1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09658__A _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16378_ clknet_leaf_62_wb_clk_i _02132_ _00361_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[101\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_42_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08562__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08082__A0 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15329_ net1240 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__inv_2
XANTENNA__11700__B net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18048_ net1548 vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__buf_2
XANTENNA__09096__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11508__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10035__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout406 _03565_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_4
X_09821_ _05491_ _06160_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__xor2_2
Xfanout417 _03562_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_8
XFILLER_0_26_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09582__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout428 _07965_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout439 _07962_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_6
XANTENNA__12023__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[20\] net806 net738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__a22o_1
XANTENNA__10332__A _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13130__B2 team_01_WB.instance_to_wrap.a1.ADR_I\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08703_ net601 net583 _05041_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_119_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12958__S net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09683_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[22\] net800 net799 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__a22o_1
XANTENNA__11862__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08634_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[10\] net901
+ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08737__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[19\] net938 vssd1
+ vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout442_A _07962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1184_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10247__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08496_ _04827_ _04828_ _04829_ _04835_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__or4_1
XFILLER_0_71_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10798__A3 _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12693__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1351_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout707_A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09568__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08472__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13736__A3 _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08903__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09117_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[14\] net894
+ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_1333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08612__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09048_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[12\] net883 vssd1
+ vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17878__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold460 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold471 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08376__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11010_ _05682_ net511 vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__nor2_1
Xhold493 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09734__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17108__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout951 _04658_ vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__buf_4
XFILLER_0_95_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout962 _04648_ vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13657__C1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout973 _04633_ vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__buf_4
XFILLER_0_95_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout984 _04499_ vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout995 net996 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09325__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12961_ net1811 net872 net359 _03715_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09876__A1 _06215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1160 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 _02088_ vssd1 vssd1 vccd1 vccd1 net2787 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ net1319 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__inv_2
X_11912_ net2168 net288 net482 vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1182 team_01_WB.instance_to_wrap.cpu.f0.num\[20\] vssd1 vssd1 vccd1 vccd1 net2798
+ sky130_fd_sc_hd__dlygate4sd3_1
X_15680_ net1238 vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__inv_2
XANTENNA__11683__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12892_ _05678_ net578 vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__nor2_1
Xhold1193 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ net1274 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ net2385 net231 net489 vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ clknet_leaf_42_wb_clk_i _03037_ _01333_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10238__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11435__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ net1388 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11774_ net2280 net263 net495 vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__mux2_1
X_16301_ clknet_leaf_75_wb_clk_i net1784 _00284_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13513_ net722 _07088_ net1067 vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__o21a_1
X_17281_ clknet_leaf_48_wb_clk_i _02968_ _01264_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10725_ _07060_ _07064_ net530 vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14493_ net1398 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16232_ clknet_leaf_106_wb_clk_i net1858 _00220_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
X_13444_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] _05419_ vssd1 vssd1
+ vccd1 vccd1 _03905_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10656_ net523 _06988_ _06991_ _06906_ net339 vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__o221a_1
XFILLER_0_36_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11738__A2 _07449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16163_ clknet_leaf_102_wb_clk_i _01926_ _00151_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11520__B net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10587_ _06883_ net337 _06916_ _06926_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__a211o_1
X_13375_ net1691 net830 _03838_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1
+ vccd1 vccd1 _01872_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12108__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10417__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15114_ net1276 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__inv_2
X_12326_ net2789 net225 net427 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__mux2_1
X_16094_ clknet_leaf_102_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[16\]
+ _00082_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11947__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15045_ net1208 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12257_ net3162 net291 net440 vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11208_ _06920_ _07050_ _07026_ vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__a21bo_1
X_12188_ net2097 net317 net449 vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__mux2_1
XANTENNA__13447__B _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11139_ net516 _06924_ vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__nor2_1
X_16996_ clknet_leaf_54_wb_clk_i _02683_ _00979_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09316__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15947_ net1403 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13463__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15878_ net1387 vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08557__A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14829_ net1212 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__inv_2
X_17617_ clknet_leaf_110_wb_clk_i _03302_ _01558_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16625__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10229__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08350_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[30\] net799 net778 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17548_ clknet_leaf_131_wb_clk_i _03235_ _01531_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08281_ net1815 net1756 net1046 vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17479_ clknet_leaf_16_wb_clk_i _03166_ _01462_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09388__A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08292__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16775__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08723__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12018__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11857__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_2
XANTENNA__09555__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout214 _07838_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_2
XANTENNA_fanout392_A _03568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout225 net226 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_2
Xfanout236 net238 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_2
X_09804_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[14\] net805 net795 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__a22o_1
Xfanout247 net250 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_2
Xfanout258 _07892_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_2
Xfanout269 net270 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_2
X_07996_ team_01_WB.instance_to_wrap.cpu.f0.num\[28\] vssd1 vssd1 vccd1 vccd1 _04494_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_66_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17400__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[20\] net946
+ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__and3_1
XANTENNA__12688__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13654__A2 _07449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1399_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10468__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09666_ net1120 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[22\] net949
+ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__and3_1
X_08617_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[11\] net696 net665 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[11\]
+ _04956_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09597_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[24\] net964
+ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08548_ net1071 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[19\] net922
+ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__and3_1
XANTENNA__11324__C team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08479_ net1083 net892 vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__and2_2
XFILLER_0_108_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10510_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[31\] net821 _06830_ _06833_
+ _06841_ vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_135_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11490_ net367 _07772_ net3279 net874 vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_80_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08633__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10441_ net504 _06780_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__nor2_1
XANTENNA__08046__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14119__B1 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13590__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13160_ net115 net843 net840 net2036 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10372_ _06708_ _06710_ _06711_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__or3_1
XANTENNA__08930__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12111_ net2125 net287 net457 vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__mux2_1
XANTENNA__11767__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13091_ _03714_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\] net861 vssd1 vssd1
+ vccd1 vccd1 _02034_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_10__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09546__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ net2862 net232 net466 vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__mux2_1
Xhold290 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16850_ clknet_leaf_135_wb_clk_i _02537_ _00833_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout770 _04672_ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__clkbuf_8
X_15801_ net1323 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__inv_2
Xfanout781 _04663_ vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_4
Xfanout792 net793 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16781_ clknet_leaf_2_wb_clk_i _02468_ _00764_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13993_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[88\] _04240_ _04243_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[24\]
+ _04284_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__a221o_1
XANTENNA__09849__A1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12598__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13645__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16648__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13283__A _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15732_ net1267 vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[9\] net1036 vssd1 vssd1 vccd1
+ vccd1 _03706_ sky130_fd_sc_hd__or2_1
XANTENNA__10459__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15663_ net1216 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12875_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[30\] _03657_ net1030 vssd1
+ vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17402_ clknet_leaf_59_wb_clk_i _03089_ _01385_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14614_ net1361 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__inv_2
XANTENNA__11408__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11826_ net575 _07945_ _07946_ vssd1 vssd1 vccd1 vccd1 _07947_ sky130_fd_sc_hd__and3_4
X_15594_ net1273 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16798__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14070__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17333_ clknet_leaf_122_wb_clk_i _03020_ _01316_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14545_ net1399 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11757_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07942_ sky130_fd_sc_hd__and2b_2
XFILLER_0_44_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10092__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17264_ clknet_leaf_126_wb_clk_i _02951_ _01247_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10708_ net336 _07045_ _07047_ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14476_ net1390 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09639__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11688_ net612 _07810_ _07887_ _07886_ vssd1 vssd1 vccd1 vccd1 _07888_ sky130_fd_sc_hd__a31o_4
XFILLER_0_70_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12908__A1 _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09001__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16215_ clknet_leaf_79_wb_clk_i _01975_ _00203_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08037__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13427_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] _04971_ vssd1 vssd1
+ vccd1 vccd1 _03888_ sky130_fd_sc_hd__xor2_1
X_10639_ net527 _06928_ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__and2_1
X_17195_ clknet_leaf_3_wb_clk_i _02882_ _01178_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13581__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16146_ clknet_leaf_96_wb_clk_i _01909_ _00134_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13358_ net585 _07686_ _03829_ _03828_ net564 vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12309_ net2938 net261 net432 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16077_ clknet_leaf_95_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_atmax _00065_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.enable sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13289_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] _03751_ vssd1 vssd1 vccd1 vccd1
+ _03776_ sky130_fd_sc_hd__or2_1
XANTENNA__16178__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13333__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15028_ net1267 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__inv_2
XANTENNA__17423__CLK clknet_leaf_143_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09671__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16979_ clknet_leaf_135_wb_clk_i _02666_ _00962_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_1
X_09520_ _05856_ _05857_ _05858_ _05859_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__or4_1
XANTENNA__17573__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12301__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08718__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09451_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[29\] net670 _05782_ _05789_
+ _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_56_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08402_ net1155 _04727_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__nand2_1
XANTENNA__10870__A2 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09382_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[26\] net939 net664 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[26\]
+ net707 vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09068__A2 _04776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14061__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08276__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08333_ net988 net941 vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout238_A _07873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10083__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08264_ net2244 net2164 net1050 vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08226__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08195_ net2589 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[78\] net1044 vssd1 vssd1
+ vccd1 vccd1 _03492_ sky130_fd_sc_hd__mux2_1
XANTENNA__09225__C1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout405_A _03565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1147_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08579__A1 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09776__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09240__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1314_A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09284__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1009 net1014 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11886__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13815__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout941_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ team_01_WB.instance_to_wrap.cpu.f0.i\[17\] vssd1 vssd1 vccd1 vccd1 _04477_
+ sky130_fd_sc_hd__inv_2
X_09718_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[21\] net740 _06037_ _06045_
+ _06047_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12211__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10990_ _07318_ _07329_ net541 vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08503__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09649_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[23\] net735 _05976_ _05978_
+ _05979_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14037__C1 _04152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12660_ net2897 net248 net389 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11611_ _07824_ _07826_ net614 vssd1 vssd1 vccd1 vccd1 _07827_ sky130_fd_sc_hd__mux2_4
XFILLER_0_33_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12591_ net2189 net222 net397 vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14330_ net1344 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11542_ net2441 net1158 net588 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] vssd1
+ vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17913__1429 vssd1 vssd1 vccd1 vccd1 _17913__1429/HI net1429 sky130_fd_sc_hd__conb_1
X_14261_ net1311 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__inv_2
X_11473_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[26\] net580 vssd1 vssd1 vccd1
+ vccd1 _07764_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_59_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16000_ net1337 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__inv_2
XANTENNA_input70_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ net27 net838 _03738_ net3095 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__a22o_1
XANTENNA__13563__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[27\] net796 _06751_ _06756_
+ _06758_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09756__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14192_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\] _04458_ net1410 vssd1
+ vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ net75 net849 net634 net1830 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10355_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[17\] net782 _06681_ _06682_
+ _06686_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_81_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09519__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13074_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[12\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[20\]
+ net854 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__mux2_1
X_17951_ net1451 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
X_10286_ _06622_ _06623_ _06624_ _06625_ vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09194__C _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16902_ clknet_leaf_41_wb_clk_i _02589_ _00885_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16470__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12025_ net575 _07942_ _07951_ vssd1 vssd1 vccd1 vccd1 _07954_ sky130_fd_sc_hd__and3_1
XANTENNA__17596__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17882_ clknet_leaf_106_wb_clk_i _03557_ _01822_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10133__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16833_ clknet_leaf_43_wb_clk_i _02520_ _00816_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09922__C net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13618__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16764_ clknet_leaf_32_wb_clk_i _02451_ _00747_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12121__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13976_ _04219_ _04220_ _04237_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__and3_4
XFILLER_0_57_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15715_ net1175 vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__inv_2
X_12927_ net1029 _03652_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__and2_2
XFILLER_0_53_1516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16695_ clknet_leaf_136_wb_clk_i _02382_ _00678_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11960__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11061__A2_N _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15646_ net1263 vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12858_ net2275 net281 net379 vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__mux2_1
XANTENNA__14043__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ net3096 net260 net493 vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15577_ net1255 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12789_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[13\] _07553_ net1028 vssd1 vssd1
+ vccd1 vccd1 _03621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17316_ clknet_leaf_53_wb_clk_i _03003_ _01299_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14528_ net1383 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17247_ clknet_leaf_24_wb_clk_i _02934_ _01230_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14459_ net1348 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09758__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13554__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10308__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09666__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17178_ clknet_leaf_58_wb_clk_i _02865_ _01161_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09222__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10907__A3 _07014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16129_ clknet_leaf_91_wb_clk_i _00020_ _00117_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08951_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[6\] net653 _05279_ _05281_
+ _05284_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_45_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08882_ _04755_ _05219_ _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09930__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16963__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13609__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12031__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12817__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10340__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09503_ net992 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[29\] net954 vssd1
+ vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14019__C1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13867__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11870__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1097_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ _05767_ _05769_ _05771_ _05773_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__or4_1
XFILLER_0_133_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08745__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14034__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09365_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] net712 net594 vssd1 vssd1
+ vccd1 vccd1 _05705_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08464__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08316_ net1147 net1150 net1153 net1152 vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_30_1346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_30 _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17469__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[22\] net926
+ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_25_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09461__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 _07900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_52 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_63 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ net1667 net2366 net1043 vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08178_ net2827 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[95\] net1047 vssd1 vssd1
+ vccd1 vccd1 _03509_ sky130_fd_sc_hd__mux2_1
XANTENNA__08480__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout891_A _04796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08957__D1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout989_A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16493__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12206__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10140_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[11\] net775 net747 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[11\]
+ _06479_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput181 net181 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
X_10071_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[7\] net944 vssd1
+ vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_34_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09921__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13830_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[23\] net831 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[23\] sky130_fd_sc_hd__and2_1
XANTENNA__11346__A team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13761_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_134_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10973_ _05301_ net373 vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11780__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15500_ net1219 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__inv_2
XANTENNA__10295__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12712_ net2514 net279 net383 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__mux2_1
X_16480_ clknet_leaf_108_wb_clk_i _02234_ _00463_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13692_ _04112_ _04113_ _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__or3_1
XANTENNA__14025__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_108_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15431_ net1301 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12643_ net2508 net253 net392 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_43_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09988__B1 _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11244__C1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15362_ net1267 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__inv_2
X_12574_ net2447 net256 net399 vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09452__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17101_ clknet_leaf_139_wb_clk_i _02788_ _01084_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14313_ net1350 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ net2307 net1158 net588 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1
+ vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__a22o_1
X_18081_ net1581 vssd1 vssd1 vccd1 vccd1 la_data_out[123] sky130_fd_sc_hd__buf_2
X_15293_ net1243 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17032_ clknet_leaf_22_wb_clk_i _02719_ _01015_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13536__A1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14244_ net1331 vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__inv_2
X_11456_ _04712_ _04753_ vssd1 vssd1 vccd1 vccd1 _07752_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08821__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10407_ _06641_ _06677_ _06745_ _06746_ _06639_ vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__o311a_1
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14175_ _04448_ _04449_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12116__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11387_ _04466_ _07715_ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13126_ net83 net847 net632 net1762 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__a22o_1
X_10338_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[17\] net978 vssd1
+ vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__and3_1
XANTENNA__16986__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_119_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11955__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17934_ team_01_WB.instance_to_wrap.cpu.LCD0.lcd_en vssd1 vssd1 vccd1 vccd1 net156
+ sky130_fd_sc_hd__clkbuf_1
X_13057_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[29\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[37\]
+ net854 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10269_ net1120 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[19\] net948
+ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__and3_1
Xfanout1340 net1341 vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__buf_2
XFILLER_0_20_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09912__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12008_ net2673 net266 net468 vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__mux2_1
Xfanout1351 net1359 vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__buf_4
X_17865_ clknet_leaf_82_wb_clk_i _03540_ _01805_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[4\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout1362 net1380 vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16216__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1373 net1379 vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__clkbuf_4
Xfanout1384 net1389 vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__buf_4
Xfanout1395 net1414 vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__buf_4
XFILLER_0_94_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16816_ clknet_leaf_129_wb_clk_i _02503_ _00799_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10160__A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17796_ clknet_leaf_65_wb_clk_i net2438 _01736_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13959_ _04219_ _04227_ _04237_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__and3_4
XFILLER_0_92_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16747_ clknet_leaf_4_wb_clk_i _02434_ _00730_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11690__S net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16678_ clknet_leaf_41_wb_clk_i _02365_ _00661_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16366__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14016__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09691__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15629_ net1213 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09979__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09150_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\] net703 _05486_ _05489_
+ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09099__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08101_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[9\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[8\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[11\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09081_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[13\] net896
+ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10038__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08032_ net1817 net567 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1
+ vccd1 vccd1 _03559_ sky130_fd_sc_hd__a22o_1
Xinput50 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
Xinput61 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput72 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
Xhold801 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold812 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold834 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12026__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold845 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[55\] vssd1 vssd1 vccd1 vccd1
+ net2461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 team_01_WB.instance_to_wrap.cpu.f0.num\[23\] vssd1 vssd1 vccd1 vccd1 net2472
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09983_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[2\] net822 net801 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__a22o_1
Xhold889 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11865__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[6\] net905 vssd1
+ vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1012_A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1501 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net3117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1512 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 net3128
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08865_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[3\] net890 vssd1
+ vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout472_A _07952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1523 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[18\] vssd1 vssd1 vccd1 vccd1
+ net3139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 _03469_ vssd1 vssd1 vccd1 vccd1 net3150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1545 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1556 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[25\] vssd1 vssd1 vccd1 vccd1
+ net3172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1567 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3183 sky130_fd_sc_hd__dlygate4sd3_1
X_08796_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[0\] net930 vssd1
+ vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__and3_1
X_17912__1428 vssd1 vssd1 vccd1 vccd1 _17912__1428/HI net1428 sky130_fd_sc_hd__conb_1
Xhold1578 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net3194 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10501__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1589 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net3205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12696__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1381_A net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout737_A _04687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13381__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10816__A2 _06065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08475__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14007__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17291__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09682__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08906__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09417_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] net712 net594 vssd1 vssd1
+ vccd1 vccd1 _05757_ sky130_fd_sc_hd__a21o_1
XANTENNA__13215__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout904_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11105__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09348_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[25\] net699 net695 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09279_ _05618_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08922__B net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11310_ _07648_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _07638_ vssd1
+ vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__mux2_1
XANTENNA__13518__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12290_ net2487 net291 net436 vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09737__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11529__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08641__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11241_ net336 _06919_ _07346_ vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14940__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11172_ _05417_ net342 _06912_ vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16239__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11775__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[6\] net809 _06457_ _06461_
+ _06462_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__a2111oi_1
X_15980_ net1394 vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14931_ net1234 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__inv_2
X_10054_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[0\] net743 _06374_ _06375_
+ _06378_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__a2111o_1
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09472__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11701__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14862_ net1282 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17650_ clknet_leaf_83_wb_clk_i _03335_ _01591_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10411__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16601_ clknet_leaf_51_wb_clk_i _02288_ _00584_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13813_ net1773 net833 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[6\]
+ sky130_fd_sc_hd__and2_1
X_17581_ clknet_leaf_72_wb_clk_i _03268_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dfxtp_1
XANTENNA__17634__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14793_ net1229 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16532_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[30\]
+ _00515_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13744_ team_01_WB.instance_to_wrap.cpu.RU0.state\[6\] net1061 net1167 vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_dhit sky130_fd_sc_hd__o21ba_1
X_10956_ _05043_ _06438_ vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08816__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16463_ clknet_leaf_134_wb_clk_i _02217_ _00446_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13675_ net1819 net568 net346 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1
+ vccd1 vccd1 _01827_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13206__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10887_ net516 _07023_ _07215_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15414_ net1201 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12626_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[27\] net213 net393 vssd1
+ vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__mux2_1
X_16394_ clknet_leaf_62_wb_clk_i _02148_ _00377_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[117\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09425__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15345_ net1291 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12557_ net3065 net224 net399 vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18064_ net1564 vssd1 vssd1 vccd1 vccd1 la_data_out[106] sky130_fd_sc_hd__buf_2
XANTENNA__13509__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ net1666 net876 _07758_ _07781_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__o22a_1
XFILLER_0_124_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17014__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15276_ net1181 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__inv_2
X_12488_ net3031 net291 net412 vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10991__A1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold108 _01981_ vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17015_ clknet_leaf_136_wb_clk_i _02702_ _00998_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08551__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09189__A1 _05528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14227_ net3091 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__clkbuf_1
Xhold119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11439_ net1065 _07676_ vssd1 vssd1 vccd1 vccd1 _07744_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14158_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[2\] vssd1 vssd1 vccd1 vccd1 _04439_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13109_ team_01_WB.instance_to_wrap.a1.curr_state\[2\] team_01_WB.instance_to_wrap.a1.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__nor2_2
XANTENNA__17164__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14089_ net149 net605 vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17917_ net1605 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XFILLER_0_59_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11299__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10602__B _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1170 _00026_ vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15681__A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08650_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[10\] net925
+ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1181 net1182 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__buf_4
X_17848_ clknet_leaf_75_wb_clk_i _03524_ _01788_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1192 net1194 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__buf_4
XANTENNA__10321__C net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08581_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[15\] net890
+ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__and3_1
X_17779_ clknet_leaf_71_wb_clk_i net2024 _01719_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[49\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_87_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09113__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09202_ net1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[17\] net938
+ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09416__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09133_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[14\] net890
+ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08624__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout220_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout318_A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10431__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09064_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[12\] net895
+ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__and3_1
XANTENNA__08234__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08015_ _04504_ team_01_WB.instance_to_wrap.cpu.f0.state\[7\] vssd1 vssd1 vccd1 vccd1
+ _04511_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10065__A _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold620 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14760__A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold631 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold653 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_A _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09966_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[3\] net797 _06288_ _06289_
+ _06294_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_25_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08917_ _05248_ _05254_ _05255_ _05256_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__or4_1
XANTENNA__16531__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09292__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[5\] net735 _06225_ _06228_
+ _06229_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1320 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1331 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1342 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2958 sky130_fd_sc_hd__dlygate4sd3_1
X_08848_ net602 _05153_ _05154_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_107_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1353 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[64\] vssd1 vssd1 vccd1 vccd1
+ net2969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2980 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1375 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1386 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3002 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13823__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1397 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3013 sky130_fd_sc_hd__dlygate4sd3_1
X_08779_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[0\] net901 vssd1
+ vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__and3_1
XANTENNA__16681__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10810_ net531 _05261_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__nand2_1
XANTENNA__11624__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11790_ net2763 net292 net496 vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08636__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10741_ _06983_ _06985_ net537 vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__mux2_1
XANTENNA__11462__A2 _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14935__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13460_ _03856_ _03858_ _03919_ _04847_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__a32o_1
X_10672_ net550 _06366_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__nor2_1
XANTENNA__17037__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09407__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12411_ net2854 net227 net420 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08615__B1 _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] _05705_ vssd1 vssd1
+ vccd1 vccd1 _03852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15130_ net1190 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12342_ net2627 net259 net430 vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15061_ net1221 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__inv_2
XANTENNA__17187__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12273_ net2416 net269 net435 vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__mux2_1
X_14012_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[89\] _04241_ _04244_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[97\]
+ _04293_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11224_ net523 _07124_ _07563_ vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09040__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10725__A1 _07064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12902__B net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09591__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ _07211_ _07214_ net517 vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10106_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[6\] net745 net734 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15963_ net1403 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11086_ _05805_ net513 vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__nor2_1
XANTENNA__13675__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17702_ clknet_leaf_101_wb_clk_i _03386_ _01643_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_10037_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[0\] net975 vssd1
+ vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14914_ net1266 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
X_15894_ net1391 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09894__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17633_ clknet_leaf_115_wb_clk_i _03318_ _01574_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\]
+ sky130_fd_sc_hd__dfrtp_4
X_14845_ net1262 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17564_ clknet_leaf_59_wb_clk_i _03251_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14776_ net1199 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11988_ net2134 net308 net474 vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__mux2_1
XANTENNA__09646__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09004__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08546__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16515_ clknet_leaf_111_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[13\]
+ _00498_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13727_ _03735_ _04098_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__nand2_1
X_10939_ _07185_ _07278_ _07276_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11453__A2 _04621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17495_ clknet_leaf_136_wb_clk_i _03182_ _01478_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10661__A0 _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16446_ clknet_leaf_44_wb_clk_i _02200_ _00429_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13658_ net187 _04089_ _04090_ net727 vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_136_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12609_ net2690 net227 net396 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16377_ clknet_leaf_65_wb_clk_i _02131_ _00360_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[100\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11205__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08606__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13589_ net199 net195 _07811_ _07883_ net645 vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_14_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15328_ net1241 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_41_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12953__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_134_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_134_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10964__B2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17911__1427 vssd1 vssd1 vccd1 vccd1 _17911__1427/HI net1427 sky130_fd_sc_hd__conb_1
X_18047_ net1547 vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__buf_2
XFILLER_0_83_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15259_ net1181 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10316__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09674__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09820_ net377 _05378_ _05416_ _05454_ _04749_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__a41o_1
Xfanout407 _03564_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_8
Xfanout418 _03562_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12304__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout429 _07965_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_8
X_09751_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[20\] _04636_ net754
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[20\] vssd1 vssd1 vccd1 vccd1
+ _06091_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08702_ net601 net583 _05041_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__a21o_1
X_09682_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[22\] net807 net788 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__a22o_1
XANTENNA__11141__A1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08542__C1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[10\] net892 vssd1
+ vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_102_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08564_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[19\] net697 _04901_
+ _04902_ _04903_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14091__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08845__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08495_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[23\] net687 _04784_ _04822_
+ net706 vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout435_A _07963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1177_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13197__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout602_A _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09116_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] _04846_ net593 vssd1 vssd1
+ vccd1 vccd1 _05456_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_21_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08073__B2 team_01_WB.instance_to_wrap.cpu.f0.write_data\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09287__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold1452_A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09047_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[12\] net927
+ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold450 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 net2066
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13818__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10707__B2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold483 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold494 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12214__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10523__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10183__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout930 net933 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_4
Xfanout941 net942 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_4
XFILLER_0_95_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09949_ net993 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[3\] net950 vssd1
+ vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__and3_1
Xfanout952 _04658_ vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__clkbuf_4
Xfanout963 _04648_ vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout974 _04633_ vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__buf_2
Xfanout985 net987 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[2\] _05258_ net1035 vssd1
+ vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout996 net1014 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1150 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2766 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ net2522 net257 net481 vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__mux2_1
Xhold1161 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2777 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1172 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2788 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12880__A1 _05779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1183 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2799 sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ net1801 net873 net360 _03668_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a22o_1
Xhold1194 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2810 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ net1228 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11354__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ net2802 net266 net489 vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__mux2_1
XANTENNA__14082__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09628__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14561_ net1402 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__inv_2
XANTENNA__11073__B _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ net1766 net270 net495 vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16427__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14665__A net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10643__A0 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16300_ clknet_leaf_79_wb_clk_i net3114 _00283_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13512_ net185 _03968_ _03969_ net725 vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__a211o_1
XFILLER_0_137_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17280_ clknet_leaf_29_wb_clk_i _02967_ _01263_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10724_ _07061_ _07063_ net519 vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09759__A _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14492_ net1390 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16231_ clknet_leaf_96_wb_clk_i net1802 _00219_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13188__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13443_ _03901_ _03903_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__and2_1
X_10655_ net533 _06994_ _06993_ _05263_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_1570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16162_ clknet_leaf_96_wb_clk_i _01925_ _00150_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13374_ net1715 net830 _03838_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1
+ vccd1 vccd1 _01873_ sky130_fd_sc_hd__a22o_1
X_10586_ net503 _06882_ net335 _06925_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__a31o_1
XANTENNA__09261__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09197__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09800__A2 _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15113_ net1229 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12325_ net2242 net192 net429 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16093_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[15\]
+ _00081_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12913__A _04881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15044_ net1239 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12256_ net2324 net315 net442 vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12699__A1 _07866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11207_ _06915_ _07369_ _07371_ net336 _07546_ vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__o221a_1
X_12187_ net3160 net320 net450 vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__mux2_1
XANTENNA__10174__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11138_ _06402_ _06403_ _07477_ vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16995_ clknet_leaf_19_wb_clk_i _02682_ _00978_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_17999__1499 vssd1 vssd1 vccd1 vccd1 _17999__1499/HI net1499 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_34_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09316__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11963__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13112__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15946_ net1390 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__inv_2
X_11069_ _07408_ _07377_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_92_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09867__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17202__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15877_ net1396 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17616_ clknet_leaf_110_wb_clk_i _03301_ _01557_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13182__C net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14828_ net1184 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14073__B1 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09619__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17547_ clknet_leaf_0_wb_clk_i _03234_ _01530_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14759_ net1327 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17352__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08280_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] net1809 net1046 vssd1 vssd1
+ vccd1 vccd1 _03407_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09669__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17478_ clknet_leaf_38_wb_clk_i _03165_ _01461_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12807__B _07308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13179__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16429_ clknet_leaf_106_wb_clk_i _02183_ _00412_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17886__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08292__B net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09252__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08358__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12034__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout204 _07858_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10343__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout215 _07838_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_2
XANTENNA__10165__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout226 _07827_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_2
X_09803_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[14\] net804 net778 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[14\]
+ _06136_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__a221o_1
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_2
Xfanout248 net250 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout259 net262 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_2
X_07995_ team_01_WB.instance_to_wrap.cpu.f0.num\[30\] vssd1 vssd1 vccd1 vccd1 _04493_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout385_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11873__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ net992 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[20\] net952 vssd1
+ vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_31_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08748__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ net1120 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[22\] net978
+ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout552_A _05151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1294_A net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08616_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[11\] net685 net671 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14064__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09596_ net992 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[24\] net970 vssd1
+ vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08547_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[19\] net897 vssd1
+ vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout817_A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08478_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[23\] net910 vssd1
+ vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08483__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09491__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12209__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10518__A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13575__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10440_ _05737_ _05759_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09243__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08046__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08597__A2 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10371_ net378 _06709_ _05566_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12110_ net3011 net255 net455 vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13090_ _03713_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\] net854 vssd1 vssd1
+ vccd1 vccd1 _02035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12041_ net2735 net264 net463 vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__mux2_1
XANTENNA__11349__A team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold280 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10253__A _05374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold291 net129 vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout760 _04674_ vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11783__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout771 _04672_ vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_4
X_15800_ net1354 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__inv_2
Xfanout782 net784 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__buf_6
XFILLER_0_79_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13992_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[80\] _04245_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_85_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16780_ clknet_leaf_116_wb_clk_i _02467_ _00763_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout793 _04652_ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15731_ net1234 vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__inv_2
X_12943_ _05373_ _07757_ _03694_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_115_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11084__A _05729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17375__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15662_ net1285 vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__inv_2
X_12874_ _05833_ net580 net361 vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17401_ clknet_leaf_46_wb_clk_i _03088_ _01384_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14613_ net1367 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__inv_2
X_11825_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\]
+ vssd1 vssd1 vccd1 vccd1 _07946_ sky130_fd_sc_hd__and2b_2
X_15593_ net1230 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
XANTENNA_output102_A net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11408__A2 _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14544_ net1384 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__inv_2
X_17332_ clknet_leaf_12_wb_clk_i _03019_ _01315_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11756_ net1971 net293 net501 vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09482__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08824__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ _05805_ net331 _07044_ net369 _07046_ vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__o221a_1
X_14475_ net1395 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__inv_2
X_17263_ clknet_leaf_141_wb_clk_i _02950_ _01246_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12119__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11687_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] _07808_ vssd1 vssd1
+ vccd1 vccd1 _07887_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16214_ clknet_leaf_61_wb_clk_i net2045 _00202_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_1
X_13426_ _03885_ _03886_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10638_ _06929_ _06969_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__or2_1
XANTENNA__08037__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09234__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17194_ clknet_leaf_10_wb_clk_i _02881_ _01177_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16145_ clknet_leaf_96_wb_clk_i _01908_ _00133_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08588__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10862__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13357_ _04483_ _07684_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10569_ _06907_ _06908_ net538 vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10395__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12308_ net2629 net232 net434 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__mux2_1
X_16076_ clknet_leaf_110_wb_clk_i _01869_ _00064_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_122_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13288_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] _03746_ _03774_ vssd1 vssd1 vccd1
+ vccd1 _03775_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_127_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15027_ net1232 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15954__A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_23_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12239_ net2213 net235 net439 vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10147__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09952__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11693__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08760__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16978_ clknet_leaf_134_wb_clk_i _02665_ _00961_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_1
XFILLER_0_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15929_ net1338 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09450_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[29\] net652 net650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__a22o_1
XANTENNA__14046__B1 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08401_ _04733_ _04739_ _04740_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__and3b_1
XFILLER_0_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17868__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09381_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[26\] net904
+ net672 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[26\] vssd1 vssd1 vccd1
+ vccd1 _05721_ sky130_fd_sc_hd__a32o_1
XFILLER_0_59_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10870__A3 _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12818__A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08332_ net989 net942 vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_99_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10706__C_N net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08263_ net2229 net2248 net1044 vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12029__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10338__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16892__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08194_ net3204 net3168 net1048 vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__mux2_1
XANTENNA__09225__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_92_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_89_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11868__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout300_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13309__C1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17248__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11169__A _07269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10073__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10138__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1307_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12699__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16272__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17398__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13384__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07978_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1 _04476_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09717_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[21\] net802 net800 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__a22o_1
X_18069__1569 vssd1 vssd1 vccd1 vccd1 _18069__1569/HI net1569 sky130_fd_sc_hd__conb_1
XFILLER_0_78_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout934_A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09648_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[23\] net746 net739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__a22o_1
XANTENNA__10310__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13831__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[25\] net820 net777 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a22o_1
XANTENNA__08925__B net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11610_ _07821_ _07825_ vssd1 vssd1 vccd1 vccd1 _07826_ sky130_fd_sc_hd__and2b_1
XANTENNA__11632__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12590_ net3231 net224 net395 vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08644__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09102__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11541_ net2840 net1159 net588 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1
+ vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10248__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17998__1498 vssd1 vssd1 vccd1 vccd1 _17998__1498/HI net1498 sky130_fd_sc_hd__conb_1
XFILLER_0_11_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14260_ net1311 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11472_ net368 _07763_ net1757 net875 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08941__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11778__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13211_ net28 net836 net629 net2585 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__o22a_1
X_10423_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[27\] net762 net752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14191_ _04458_ _04459_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__nor2_1
XANTENNA__13563__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10682__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13142_ net86 net849 net634 net1753 vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input63_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[17\] net760 _06680_
+ _06684_ _06690_ vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09475__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13073_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[21\]
+ net854 vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__mux2_1
X_17950_ net1450 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XANTENNA__16615__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10285_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[19\] net791 net750 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__a22o_1
XANTENNA__10414__C net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11326__B2 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16901_ clknet_leaf_39_wb_clk_i _02588_ _00884_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12024_ net3183 net292 net468 vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17881_ clknet_leaf_104_wb_clk_i _03556_ _01821_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_16832_ clknet_leaf_29_wb_clk_i _02519_ _00815_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_137_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12402__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 _07785_ vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16765__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08819__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16763_ clknet_leaf_50_wb_clk_i _02450_ _00746_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12826__A1 _07489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13975_ _04217_ _04219_ _04227_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__and3_4
XFILLER_0_87_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15714_ net1265 vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12926_ net2636 net870 net357 _03693_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a22o_1
X_16694_ clknet_leaf_1_wb_clk_i _02381_ _00677_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15645_ net1250 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__inv_2
X_12857_ net3151 net302 net382 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11808_ net2470 net233 net492 vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15576_ net1183 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__inv_2
X_12788_ net2261 net641 net608 _03620_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09012__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11262__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17315_ clknet_leaf_19_wb_clk_i _03002_ _01298_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08554__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14527_ net1332 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11739_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\]
+ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1 vccd1 vccd1 _07929_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17246_ clknet_leaf_48_wb_clk_i _02933_ _01229_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09947__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16145__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08851__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14458_ net1348 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13409_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] _05220_ vssd1 vssd1 vccd1
+ vccd1 _03870_ sky130_fd_sc_hd__and2_1
XANTENNA__13554__A2 _07621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13469__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17177_ clknet_leaf_58_wb_clk_i _02864_ _01160_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14389_ net1304 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16128_ clknet_leaf_91_wb_clk_i _00019_ _00116_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16295__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08950_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[6\] net661 _05272_ _05273_
+ _05289_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_121_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16059_ clknet_leaf_89_wb_clk_i _01852_ _00047_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10324__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08881_ net602 _05220_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12312__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17690__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09502_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[29\] net971
+ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10828__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08497__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14019__B1 _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[28\] net693 net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[28\]
+ _05772_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout250_A _07842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09364_ _05691_ _05692_ _05703_ net704 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__o32a_4
XANTENNA__13242__B2 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11171__B _06924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08315_ net1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[30\] net957
+ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12982__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_20 _07827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[22\] net922
+ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_31 _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout515_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1257_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_42 _07900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[35\] net3166 net1051 vssd1 vssd1
+ vccd1 vccd1 _03441_ sky130_fd_sc_hd__mux2_1
XANTENNA__09857__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_64 _07566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17070__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08177_ net2542 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[96\] net1042 vssd1 vssd1
+ vccd1 vccd1 _03510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10359__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12753__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09295__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
XFILLER_0_80_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput182 net182 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XANTENNA__09592__A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ _06406_ _06408_ _06254_ _06285_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__o211ai_4
XANTENNA__13826__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08724__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__C1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12222__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10531__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08639__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11346__B team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13744__B1_N net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08001__A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13760_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_74_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10972_ _05301_ net373 vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__or2_1
XANTENNA__13481__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09685__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10295__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12711_ net3228 net302 net384 vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__mux2_1
XANTENNA__11492__B1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13691_ team_01_WB.instance_to_wrap.cpu.c0.count\[11\] team_01_WB.instance_to_wrap.cpu.c0.count\[8\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[7\] team_01_WB.instance_to_wrap.cpu.c0.count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_78_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15430_ net1324 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__inv_2
X_12642_ net2640 net227 net392 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09437__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17413__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15361_ net1247 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__inv_2
X_12573_ net2570 net260 net400 vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__mux2_1
X_17100_ clknet_leaf_131_wb_clk_i _02787_ _01083_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11524_ net1731 net1158 net588 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1
+ vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__a22o_1
X_14312_ net1353 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18080_ net1580 vssd1 vssd1 vccd1 vccd1 la_data_out[122] sky130_fd_sc_hd__buf_2
X_15292_ net1171 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08671__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14243_ net1331 vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__inv_2
XANTENNA__13289__A team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17031_ clknet_leaf_123_wb_clk_i _02718_ _01014_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13536__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11455_ net1161 team_01_WB.instance_to_wrap.cpu.DM0.state\[2\] vssd1 vssd1 vccd1
+ vccd1 team_01_WB.instance_to_wrap.cpu.DM0.next_enable sky130_fd_sc_hd__and2_2
XFILLER_0_80_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17563__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10406_ net505 _06638_ _06675_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__o21bai_1
X_14174_ net1737 _04447_ net1169 vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11386_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] net1062 _07668_ _07714_ vssd1
+ vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__nand4_2
XFILLER_0_110_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13125_ net84 net847 net632 net1865 vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10337_ _06675_ _06676_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13056_ net2656 net1673 net852 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__mux2_1
X_17933_ net1435 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
X_10268_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[19\] net802 _06605_
+ _06606_ _06607_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__a2111o_1
Xfanout1330 net1331 vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__buf_4
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12007_ net2002 net268 net467 vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__mux2_1
Xfanout1341 net1342 vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17864_ clknet_leaf_81_wb_clk_i _03539_ _01804_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10441__A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12132__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1352 net1358 vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__buf_4
X_10199_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[8\] net953 vssd1
+ vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__and3_1
Xfanout1363 net1380 vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__buf_4
Xfanout1374 net1375 vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__buf_4
Xfanout1385 net1389 vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__buf_4
X_16815_ clknet_leaf_143_wb_clk_i _02502_ _00798_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1396 net1404 vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__buf_4
X_17795_ clknet_leaf_69_wb_clk_i net2069 _01735_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11971__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16746_ clknet_leaf_11_wb_clk_i _02433_ _00729_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13958_ _04238_ _04248_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__nor2_4
XFILLER_0_88_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09676__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09441__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09140__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12909_ net2308 net870 net357 _03681_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a22o_1
X_16677_ clknet_leaf_31_wb_clk_i _02364_ _00660_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13889_ net1329 _04146_ _04195_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__nor3_1
XFILLER_0_115_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15628_ net1220 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__inv_2
XANTENNA__09428__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13224__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15559_ net1300 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08100_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[3\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[2\]
+ _04569_ _04570_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__or4_1
X_09080_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[13\] net902
+ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08031_ net1747 net567 net346 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1
+ vccd1 vccd1 _03560_ sky130_fd_sc_hd__a22o_1
Xinput40 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_2
X_17229_ clknet_leaf_138_wb_clk_i _02916_ _01212_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12307__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18068__1568 vssd1 vssd1 vccd1 vccd1 _18068__1568/HI net1568 sky130_fd_sc_hd__conb_1
Xinput51 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_1
Xhold802 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
Xinput62 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11538__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xinput73 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_1
Xhold813 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[8\] vssd1 vssd1 vccd1 vccd1
+ net2429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09600__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold835 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 _02094_ vssd1 vssd1 vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08954__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09982_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[2\] net792 net777 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold868 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold879 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08933_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[6\] net908 vssd1
+ vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout298_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13160__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08864_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[3\] net932 vssd1
+ vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__and3_1
Xhold1502 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3118 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12042__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1513 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net3129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1524 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[65\] vssd1 vssd1 vccd1 vccd1
+ net3140 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1005_A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1535 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3151 sky130_fd_sc_hd__dlygate4sd3_1
X_17997__1497 vssd1 vssd1 vccd1 vccd1 _17997__1497/HI net1497 sky130_fd_sc_hd__conb_1
Xhold1546 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1557 _02064_ vssd1 vssd1 vccd1 vccd1 net3173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08795_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[0\] net909 vssd1
+ vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__and3_1
Xhold1568 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net3184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1579 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3195 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11881__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout465_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08756__A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16310__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10816__A3 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout632_A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08475__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\] net704 _05749_ _05755_
+ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__o22a_2
XFILLER_0_109_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13215__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15589__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09347_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[25\] net688 net686 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13620__D1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09278_ net598 _05615_ _05617_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08229_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[52\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[44\]
+ net1041 vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__mux2_1
XANTENNA__13518__A2 _07566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12217__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11529__B2 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11240_ _06750_ _06817_ _06822_ net344 vssd1 vssd1 vccd1 vccd1 _07580_ sky130_fd_sc_hd__a31o_1
X_11171_ _05416_ _06924_ vssd1 vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10122_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[6\] net777 net749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__a22o_1
XANTENNA__13151__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14930_ net1232 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10053_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[0\] net821 net795 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__a22o_1
XANTENNA__10504__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11701__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ net1210 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ clknet_leaf_27_wb_clk_i _02287_ _00583_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13812_ net2901 net833 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[5\]
+ sky130_fd_sc_hd__and2_1
X_17580_ clknet_leaf_71_wb_clk_i _03267_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14792_ net1276 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16531_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[29\]
+ _00514_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10955_ _05043_ _06438_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__nor2_1
X_13743_ _04136_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11092__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16803__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16462_ clknet_leaf_18_wb_clk_i _02216_ _00445_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10886_ net329 _07219_ _07221_ _07225_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__a211o_1
X_13674_ net1662 net567 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1
+ vccd1 vccd1 _01828_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15413_ net1223 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__inv_2
XANTENNA__15499__A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12625_ net1973 net218 net391 vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__mux2_1
X_16393_ clknet_leaf_65_wb_clk_i _02147_ _00376_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[116\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_109_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12965__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09497__A _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15344_ net1270 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__inv_2
X_12556_ net3008 net192 net401 vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16953__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08832__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11507_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[9\] _07756_ vssd1 vssd1 vccd1
+ vccd1 _07781_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18063_ net1563 vssd1 vssd1 vccd1 vccd1 la_data_out[105] sky130_fd_sc_hd__buf_2
XFILLER_0_53_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15275_ net1298 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__inv_2
X_12487_ net2095 net314 net414 vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12127__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17014_ clknet_leaf_140_wb_clk_i _02701_ _00997_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold109 net80 vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14226_ net3068 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__clkbuf_1
X_11438_ _07736_ _07743_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11966__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14157_ _04195_ _04438_ net1411 vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17309__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11369_ _07670_ _07697_ vssd1 vssd1 vccd1 vccd1 _07698_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13108_ team_01_WB.EN_VAL_REG net72 _03730_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__mux2_1
X_14088_ _04348_ _04375_ _04356_ net1169 vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__o211a_1
XANTENNA__13466__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09663__C net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13142__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17916_ net1604 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15962__A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13039_ net2663 net2461 net861 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1160 team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1 net1160
+ sky130_fd_sc_hd__buf_2
XANTENNA__17459__CLK clknet_leaf_137_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1171 net1173 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__buf_4
XANTENNA__09361__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17847_ clknet_leaf_63_wb_clk_i _03523_ _01787_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[117\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1182 net1185 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__clkbuf_2
Xfanout1193 net1194 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__buf_2
XFILLER_0_117_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08580_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[15\] net681 net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__a22o_1
X_17778_ clknet_leaf_76_wb_clk_i _03454_ _01718_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09113__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16729_ clknet_leaf_47_wb_clk_i _02416_ _00712_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17889__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16483__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09201_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[17\] net926
+ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_100_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12956__A0 team_01_WB.instance_to_wrap.cpu.f0.write_data\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09132_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[14\] net923 vssd1
+ vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08742__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09063_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[12\] _04767_
+ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__and3_1
XANTENNA__12037__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10346__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08014_ team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] vssd1 vssd1 vccd1 vccd1 _04510_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_13_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold610 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold621 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold632 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[10\] vssd1 vssd1 vccd1 vccd1
+ net2248 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11876__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold643 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold654 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold665 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1122_A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold676 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold687 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[72\] vssd1 vssd1 vccd1 vccd1
+ net2303 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08250__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold698 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[3\] net823 _06287_ _06290_
+ _06296_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09573__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13133__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[2\] net674 _05226_ _05228_
+ _05233_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__a2111o_1
X_09896_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[5\] net808 _06223_ _06224_
+ _06231_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__a2111o_1
Xhold1310 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1321 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1332 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2948 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09352__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ _05178_ _05182_ _05186_ _05155_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__o31a_4
Xhold1343 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1354 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[118\] vssd1 vssd1 vccd1 vccd1
+ net2970 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout847_A net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13392__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1365 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1376 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2992 sky130_fd_sc_hd__dlygate4sd3_1
X_08778_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[0\] net913 vssd1
+ vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__and3_1
XANTENNA__12500__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1387 team_01_WB.instance_to_wrap.cpu.f0.num\[6\] vssd1 vssd1 vccd1 vccd1 net3003
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1398 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3014 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09104__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11447__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13987__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10740_ _06982_ _06999_ net533 vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16976__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10671_ _07010_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12410_ net2507 net289 net421 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__mux2_1
XANTENNA__11640__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13390_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] _05705_ vssd1 vssd1
+ vccd1 vccd1 _03851_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09812__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10958__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08652__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14149__C1 _04152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12341_ net2126 net232 net429 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15060_ net1267 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__inv_2
X_12272_ net2927 net237 net435 vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__mux2_1
X_14011_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[41\] _04246_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[113\]
+ _04292_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__a221o_1
XANTENNA__11786__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08918__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ _06890_ _06906_ _06909_ _05263_ net339 vssd1 vssd1 vccd1 vccd1 _07563_ sky130_fd_sc_hd__o221a_1
XFILLER_0_31_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10186__B1 _06502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11922__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16356__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08160__S net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ net345 _07492_ _07493_ vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__or3_1
XANTENNA__09591__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13124__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10105_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[6\] net823 net797 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[6\]
+ _06443_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__a221o_1
X_15962_ net1391 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__inv_2
X_11085_ _05759_ net504 _07347_ _07423_ _07424_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__o221a_1
XANTENNA__13675__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17701_ clknet_leaf_101_wb_clk_i _03385_ _01642_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10422__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[0\] net943 vssd1
+ vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__and3_1
X_14913_ net1246 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__inv_2
XANTENNA__11686__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15893_ net1406 vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ clknet_leaf_117_wb_clk_i _03317_ _01573_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12410__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14844_ net1171 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18067__1567 vssd1 vssd1 vccd1 vccd1 _18067__1567/HI net1567 sky130_fd_sc_hd__conb_1
XFILLER_0_86_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08827__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17563_ clknet_leaf_60_wb_clk_i _03250_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13978__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08839__D1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14775_ net1199 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__inv_2
X_11987_ net2216 net312 net472 vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16514_ clknet_leaf_111_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[12\]
+ _00497_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13726_ team_01_WB.instance_to_wrap.cpu.DM0.dhit net2220 _04575_ vssd1 vssd1 vccd1
+ vccd1 _00018_ sky130_fd_sc_hd__a21o_1
XANTENNA__10110__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10938_ net526 _07277_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17494_ clknet_leaf_141_wb_clk_i _03181_ _01477_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10661__A1 _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16445_ clknet_leaf_33_wb_clk_i _02199_ _00428_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13657_ net199 net195 _07934_ net645 vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__o211a_1
X_10869_ _06715_ _06740_ _07112_ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__nand3_2
XFILLER_0_67_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12608_ net2142 net288 net397 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08606__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16376_ clknet_leaf_73_wb_clk_i net2384 _00359_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09803__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13588_ _03901_ _04032_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09020__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18115_ net637 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_41_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08562__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15327_ net1256 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_41_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12539_ net2651 net231 net406 vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__mux2_1
X_17996__1496 vssd1 vssd1 vccd1 vccd1 _17996__1496/HI net1496 sky130_fd_sc_hd__conb_1
XANTENNA__14861__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18046_ net1546 vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__buf_2
XANTENNA__14155__A2 _04195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09955__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15258_ net1187 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08909__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14209_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] vssd1 vssd1 vccd1
+ vccd1 _02278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15189_ net1220 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17281__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout408 _03564_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_4
XANTENNA__09582__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout419 net422 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_103_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13115__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09750_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[20\] net808 net796 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__a22o_1
XANTENNA__11126__C1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09334__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08701_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] net596 net601 vssd1 vssd1
+ vccd1 vccd1 _05041_ sky130_fd_sc_hd__a21oi_1
X_09681_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[22\] net821 net768 _06011_
+ _06014_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_94_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08542__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[10\] net906
+ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__and3_1
XANTENNA__12320__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08737__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16999__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08563_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[19\] net882
+ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__and3_1
XANTENNA__11444__B net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08494_ _04830_ _04831_ _04832_ _04833_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16229__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout428_A _07965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09568__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09115_ _05454_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__inv_2
XANTENNA__08472__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10404__A1 _06598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14771__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10076__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1337_A net1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16379__CLK clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09046_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[12\] net891
+ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13387__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold440 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10804__A _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold451 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09076__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold462 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 net2078
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10707__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold473 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold495 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[20\] vssd1 vssd1 vccd1 vccd1
+ net2111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout964_A _04645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout920 net921 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_4
Xfanout931 net933 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09948_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[3\] _04665_
+ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__and3_1
Xfanout942 _04671_ vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13657__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout953 net954 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_8
Xfanout964 _04645_ vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__buf_4
Xfanout975 _04631_ vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__buf_4
Xfanout986 net987 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09325__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _06216_ _06217_ vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout997 net999 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2767 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ net3256 net261 net482 vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2778 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12230__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1173 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2789 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[25\] _03667_ net1032 vssd1
+ vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__mux2_1
XANTENNA__17004__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1184 team_01_WB.instance_to_wrap.cpu.c0.count\[8\] vssd1 vssd1 vccd1 vccd1 net2800
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1195 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2811 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08647__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10891__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ net2081 net267 net487 vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14560_ net1383 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11772_ net2187 net237 net495 vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08944__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10723_ _07062_ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10643__A1 _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13511_ net197 net193 _07834_ net643 vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_1362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14491_ net1407 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_109_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16230_ clknet_leaf_105_wb_clk_i _01990_ _00218_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13442_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] _05456_ vssd1 vssd1
+ vccd1 vccd1 _03903_ sky130_fd_sc_hd__xnor2_1
X_10654_ _05898_ net504 net543 vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16161_ clknet_leaf_102_wb_clk_i _01924_ _00149_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13373_ net2072 net830 _03838_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1
+ vccd1 vccd1 _01874_ sky130_fd_sc_hd__a22o_1
X_10585_ _06882_ net332 _06922_ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15112_ net1287 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__inv_2
XANTENNA__10417__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12324_ _07790_ _07794_ net573 vssd1 vssd1 vccd1 vccd1 _07965_ sky130_fd_sc_hd__and3_4
XFILLER_0_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_1_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16092_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[14\]
+ _00080_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12255_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[2\] net320 net442 vssd1
+ vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15043_ net1188 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10159__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12405__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10714__A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11206_ _05455_ _07545_ vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12186_ net2803 net307 net450 vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_118_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ _06402_ _06403_ net345 vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_125_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16994_ clknet_leaf_35_wb_clk_i _02681_ _00977_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13648__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09316__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15945_ net1333 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__inv_2
X_11068_ _05338_ _06562_ _07259_ net340 _05374_ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_121_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[1\] net787 net734 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[1\]
+ _06344_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12140__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15876_ net1386 vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10331__B1 _06669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09015__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17615_ clknet_leaf_110_wb_clk_i _03300_ _01556_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08557__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14827_ net1297 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17546_ clknet_leaf_10_wb_clk_i _03233_ _01529_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14758_ net1325 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_127_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08854__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13709_ _04100_ _04124_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[1\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_28_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17477_ clknet_leaf_37_wb_clk_i _03164_ _01460_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14689_ net1361 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16428_ clknet_leaf_106_wb_clk_i _02182_ _00411_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_82_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16521__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16359_ clknet_leaf_67_wb_clk_i net2609 _00342_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09252__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10398__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14128__A2 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18029_ net1529 vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__buf_2
XFILLER_0_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12315__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_136_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09555__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout205 net206 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout216 _07835_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_2
X_09802_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[14\] net757 net755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[14\]
+ _06137_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout227 _07900_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_2
Xfanout238 _07873_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout249 net250 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_2
X_07994_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1 _04492_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17027__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09307__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09733_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[20\] net780 net752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout280_A _07917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11455__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_A _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12050__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ net1120 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[22\] net966
+ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__and3_1
XANTENNA__08467__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08615_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[11\] net690 _04789_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[11\] _04953_ vssd1 vssd1 vccd1
+ vccd1 _04955_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09595_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[24\] net822 net799 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_71_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout545_A _05152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1287_A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08546_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[19\] net931 vssd1
+ vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08477_ net1004 net909 vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout712_A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08483__B net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09298__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire617 _05335_ vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15597__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08046__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14119__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10370_ net378 _05566_ _06709_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13829__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08930__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09029_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[9\] net661 _05346_ _05356_
+ _05357_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_32_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18066__1566 vssd1 vssd1 vccd1 vccd1 _18066__1566/HI net1566 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_72_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10421__A_N net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12040_ net2021 net268 net463 vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__mux2_1
Xhold270 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[24\] vssd1 vssd1 vccd1 vccd1 net1886
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09546__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold281 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _01995_ vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12550__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_127_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout750 _04680_ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08939__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout761 _04674_ vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout772 net774 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_6
Xfanout783 net784 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__buf_6
X_13991_ _04279_ _04280_ _04281_ _04282_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__or4_1
Xfanout794 net797 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15730_ net1233 vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12942_ net359 _03703_ _03704_ net872 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a32o_1
X_17995__1495 vssd1 vssd1 vccd1 vccd1 _17995__1495/HI net1495 sky130_fd_sc_hd__conb_1
XFILLER_0_73_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11084__B _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15661_ net1211 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__inv_2
X_12873_ net2001 net870 net357 _03656_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__a22o_1
X_17400_ clknet_leaf_30_wb_clk_i _03087_ _01383_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14612_ net1365 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__inv_2
X_11824_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07945_ sky130_fd_sc_hd__and2_2
XFILLER_0_115_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15592_ net1287 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XANTENNA__08674__A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17331_ clknet_leaf_129_wb_clk_i _03018_ _01314_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14543_ net1334 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__inv_2
X_11755_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _07940_ net616 vssd1
+ vssd1 vccd1 vccd1 _07941_ sky130_fd_sc_hd__mux2_8
XANTENNA__09482__A1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11077__A_N net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17262_ clknet_leaf_8_wb_clk_i _02949_ _01245_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10706_ _05805_ _06919_ net513 vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__or3b_1
XANTENNA__10092__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14474_ net1385 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11686_ net720 _07188_ net616 _07885_ vssd1 vssd1 vccd1 vccd1 _07886_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16213_ clknet_leaf_95_wb_clk_i net1804 _00201_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13425_ _04949_ _03884_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1
+ vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__o21a_1
XANTENNA__09001__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10637_ _05835_ net331 _06976_ net369 vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__o211a_1
X_17193_ clknet_leaf_23_wb_clk_i _02880_ _01176_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16694__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16144_ clknet_leaf_96_wb_clk_i _01907_ _00132_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13356_ _07677_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10568_ net504 _06811_ net543 vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12307_ net2427 net263 net432 vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__mux2_1
X_16075_ clknet_leaf_111_wb_clk_i _01868_ _00063_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12135__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10499_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\] _04665_
+ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__and3b_1
X_13287_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] _03746_ _04518_ vssd1 vssd1 vccd1
+ vccd1 _03774_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10444__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15026_ net1233 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12238_ net3226 net239 net439 vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11974__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10552__A0 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ net2948 net272 net448 vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09671__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16977_ clknet_leaf_18_wb_clk_i _02664_ _00960_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15970__A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_15928_ net1330 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__inv_2
XANTENNA__10304__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15859_ net1396 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08400_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] _04727_ vssd1 vssd1 vccd1
+ vccd1 _04740_ sky130_fd_sc_hd__nand2_1
X_09380_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[26\] net654 net651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[26\]
+ _05719_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08584__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12818__B _07449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08331_ net1147 net1148 net1152 net1154 vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__nor4_1
X_17529_ clknet_leaf_58_wb_clk_i _03216_ _01512_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08262_ net3050 net2758 net1051 vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10083__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08193_ net1686 net2646 net1037 vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__mux2_1
XANTENNA__09225__A1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09776__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12780__A1 _07541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12045__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1035_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11169__B _07290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11335__A2 team_01_WB.instance_to_wrap.cpu.f0.state\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout495_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11884__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1202_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1 vccd1 vccd1 _04475_
+ sky130_fd_sc_hd__inv_2
X_09716_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[21\] net821 net775 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09647_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[23\] net802 net756 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14037__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09578_ _05915_ _05916_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__or3_1
XFILLER_0_72_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08529_ net1071 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[18\] net897
+ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__and3_1
XANTENNA__11632__B net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11540_ net1754 net1158 net588 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1
+ vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11471_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[27\] net580 vssd1 vssd1 vccd1
+ vccd1 _07763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13210_ net29 net838 _03738_ net2901 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a22o_1
X_10422_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\] net958
+ vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14190_ net2107 _04457_ net1169 vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12771__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13141_ net97 net850 net633 net3247 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a22o_1
X_10353_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[17\] net807 _06679_
+ _06685_ _06689_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_104_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13072_ net2234 net1625 net853 vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__mux2_1
XANTENNA__09519__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input56_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[19\] net779 net768 vssd1
+ vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__a21o_1
X_12023_ net3027 net316 net469 vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__mux2_1
X_16900_ clknet_leaf_51_wb_clk_i _02587_ _00883_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11794__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17342__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17880_ clknet_leaf_101_wb_clk_i _03555_ _01820_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10534__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16831_ clknet_leaf_7_wb_clk_i _02518_ _00814_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout580 _07752_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__buf_4
X_16762_ clknet_leaf_58_wb_clk_i _02449_ _00745_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13974_ _04217_ _04227_ _04239_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__and3_4
XFILLER_0_92_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17492__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15713_ net1246 vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__inv_2
X_12925_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[15\] _03692_ net1032 vssd1
+ vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__mux2_1
X_16693_ clknet_leaf_125_wb_clk_i _02380_ _00676_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15644_ net1173 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__inv_2
X_12856_ net2129 net285 net381 vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11807_ net1959 net264 net493 vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15575_ net1198 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12787_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] net1056 net365 _03619_
+ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17314_ clknet_leaf_34_wb_clk_i _03001_ _01297_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14526_ net1335 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11738_ net718 _07449_ net613 vssd1 vssd1 vccd1 vccd1 _07928_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11969__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17245_ clknet_leaf_40_wb_clk_i _02932_ _01228_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14457_ net1348 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11669_ _07871_ _07872_ net611 vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__mux2_2
XFILLER_0_29_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13408_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] _05112_ vssd1 vssd1 vccd1
+ vccd1 _03869_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17176_ clknet_leaf_28_wb_clk_i _02863_ _01159_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14388_ net1304 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__inv_2
XANTENNA__09666__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap714 _04726_ vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__buf_1
XFILLER_0_49_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12762__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08570__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16127_ clknet_leaf_93_wb_clk_i _00018_ _00115_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13339_ net1690 _03814_ net826 vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16058_ clknet_leaf_90_wb_clk_i _01851_ _00046_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15009_ net1247 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08880_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] net730 _05111_ net1108 vssd1
+ vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__a22o_1
XANTENNA__09930__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12817__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10340__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[29\] net946
+ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08497__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11733__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18065__1565 vssd1 vssd1 vccd1 vccd1 _18065__1565/HI net1565 sky130_fd_sc_hd__conb_1
X_09432_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[28\] net699 net675 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08745__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09203__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09363_ _05693_ _05696_ _05700_ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__or4_1
XANTENNA__10349__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout243_A _07862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08314_ net1132 net957 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__and2_2
XANTENNA__09997__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09294_ net1073 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[22\] net907
+ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_10 _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _07858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_32 _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08245_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[36\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[28\]
+ net1041 vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11879__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 _07900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout410_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1152_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_65 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout508_A _06065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08176_ net1680 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[97\] net1052 vssd1 vssd1
+ vccd1 vccd1 _03511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08480__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17994__1494 vssd1 vssd1 vccd1 vccd1 _17994__1494/HI net1494 sky130_fd_sc_hd__conb_1
XANTENNA__10764__A0 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_0_30_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout877_A team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13395__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput172 net172 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
Xoutput183 net183 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
XANTENNA__12503__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09921__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10971_ _06920_ _07141_ _07151_ _06928_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__a22o_1
XANTENNA__08488__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12710_ net3079 net286 net385 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13690_ team_01_WB.instance_to_wrap.cpu.c0.count\[14\] team_01_WB.instance_to_wrap.cpu.c0.count\[13\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[12\] team_01_WB.instance_to_wrap.cpu.c0.count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__or4b_1
XFILLER_0_6_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12641_ net2890 net288 net393 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10047__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15360_ net1243 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__inv_2
XANTENNA__09988__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11244__B2 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ net2696 net233 net402 vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11789__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14311_ net1357 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11523_ net1978 net1158 net588 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1
+ vccd1 vccd1 _03329_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15291_ net1180 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08660__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17708__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17030_ clknet_leaf_42_wb_clk_i _02717_ _01013_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14242_ net1331 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__inv_2
X_11454_ _07671_ net327 _07751_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__and3b_1
XFILLER_0_46_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10706__B _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12744__A1 _07566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10405_ _06713_ _06740_ _06712_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__o21a_1
X_14173_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[8\] _04447_ vssd1 vssd1 vccd1
+ vccd1 _04448_ sky130_fd_sc_hd__and2_1
X_11385_ _04471_ _07713_ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__nor2_2
XFILLER_0_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13124_ net1738 net847 net632 team_01_WB.instance_to_wrap.a1.ADR_I\[19\] vssd1 vssd1
+ vccd1 vccd1 _02017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10336_ _06672_ _06673_ _06674_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__nand3_1
XANTENNA__16732__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12413__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13055_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[31\] net2345 net861 vssd1 vssd1
+ vccd1 vccd1 _02070_ sky130_fd_sc_hd__mux2_1
X_17932_ net1434 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_24_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10267_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[19\] net943 vssd1
+ vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__and3_1
Xfanout1320 net1322 vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__clkbuf_4
X_12006_ net2283 net236 net467 vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__mux2_1
Xfanout1331 net1340 vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__buf_4
X_17863_ clknet_leaf_82_wb_clk_i _03538_ _01803_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[2\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout1342 net1415 vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__buf_4
X_10198_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[8\] net967 vssd1
+ vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1353 net1358 vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__buf_2
Xfanout1364 net1380 vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__buf_4
Xfanout1375 net1378 vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16882__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16814_ clknet_leaf_5_wb_clk_i _02501_ _00797_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_17794_ clknet_leaf_85_wb_clk_i _03470_ _01734_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[64\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1386 net1389 vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__buf_4
XFILLER_0_75_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1397 net1404 vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__buf_2
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16745_ clknet_leaf_9_wb_clk_i _02432_ _00728_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13957_ _04225_ _04248_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__nor2_4
XFILLER_0_53_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12908_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[20\] _03680_ net1030 vssd1
+ vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__mux2_1
X_16676_ clknet_leaf_51_wb_clk_i _02363_ _00659_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13888_ _04189_ _04194_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__nand2_4
XFILLER_0_75_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17238__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_128_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15627_ net1298 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__inv_2
X_12839_ net3017 net247 net380 vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11235__A1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09979__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15558_ net1292 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__inv_2
XANTENNA__11235__B2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08862__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11699__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14509_ net1405 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__inv_2
XANTENNA__16262__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17388__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15489_ net1249 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__inv_2
X_08030_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid _04523_ _04525_ vssd1 vssd1 vccd1
+ vccd1 _04526_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17228_ clknet_leaf_134_wb_clk_i _02915_ _01211_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput41 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput52 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12735__A1 _07019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput63 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold803 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[107\] vssd1 vssd1 vccd1 vccd1
+ net2419 sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 wbs_we_i vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
X_17159_ clknet_leaf_16_wb_clk_i _02846_ _01142_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold814 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[11\] vssd1 vssd1 vccd1 vccd1
+ net2441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold836 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[2\] net820 net783 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold869 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08932_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[6\] _04759_
+ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__and3_1
XANTENNA__11728__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12323__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09364__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08863_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[3\] net898 vssd1
+ vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__and3_1
Xhold1503 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1514 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3130 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout193_A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1525 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1536 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1547 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3163 sky130_fd_sc_hd__dlygate4sd3_1
X_08794_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[0\] net930 vssd1
+ vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__and3_1
Xhold1558 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09116__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1569 team_01_WB.instance_to_wrap.a1.BUSY_O vssd1 vssd1 vccd1 vccd1 net3185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout458_A _07956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09415_ _05751_ _05752_ _05753_ _05754_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__or4_1
XANTENNA__10079__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16605__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13215__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1367_A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09346_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[25\] net693 net676 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold1475_A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ net600 _05616_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08228_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[53\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[45\]
+ net1040 vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11529__A2 team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout994_A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08159_ net2349 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[114\] net1042 vssd1 vssd1
+ vccd1 vccd1 _03528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11170_ _06220_ _07172_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__nand2_1
XANTENNA__13837__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10121_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[6\] net801 _06458_ _06460_
+ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__a211o_1
XFILLER_0_105_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11638__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12233__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09355__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[0\] net731 _06371_ _06372_
+ _06376_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08012__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11162__B1 _07042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11701__A2 _07207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14860_ net1209 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
XANTENNA__08947__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16135__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14100__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13811_ net2585 net834 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[4\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_19_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14791_ net1327 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__inv_2
XANTENNA__10688__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16530_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[28\]
+ _00513_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11373__A team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13742_ net1160 net1026 vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__and2b_1
XANTENNA__10268__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08158__S net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ _07292_ _07293_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__xor2_1
XFILLER_0_54_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16461_ clknet_leaf_128_wb_clk_i _02215_ _00444_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16285__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13673_ net1669 net567 net346 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1
+ vccd1 vccd1 _01829_ sky130_fd_sc_hd__a22o_1
X_10885_ net514 _07041_ _07099_ _07224_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__a31o_1
XANTENNA__13206__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17530__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15412_ net1287 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12624_ net2291 net221 net393 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__mux2_1
X_16392_ clknet_leaf_73_wb_clk_i net3058 _00375_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15343_ net1216 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12555_ _07942_ _07951_ net574 vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__and3_4
XANTENNA__12408__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18062_ net1562 vssd1 vssd1 vccd1 vccd1 la_data_out[104] sky130_fd_sc_hd__buf_2
X_11506_ net1702 net877 _07758_ _07780_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__o22a_1
X_15274_ net1226 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12486_ net2480 net318 net414 vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17013_ clknet_leaf_126_wb_clk_i _02700_ _00996_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17680__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14225_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] vssd1 vssd1 vccd1
+ vccd1 _02262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11437_ net3245 _07700_ net326 vssd1 vssd1 vccd1 vccd1 _07743_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08397__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14156_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18064__1564 vssd1 vssd1 vccd1 vccd1 _18064__1564/HI net1564 sky130_fd_sc_hd__conb_1
XFILLER_0_21_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11368_ _07696_ vssd1 vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13107_ net73 net71 net74 _03729_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__and4_1
XANTENNA__12143__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10319_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[18\] net788 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[18\]
+ _06658_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14087_ _04365_ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__or2_2
X_11299_ net198 net194 net644 vssd1 vssd1 vccd1 vccd1 _07639_ sky130_fd_sc_hd__o21ai_2
XANTENNA__13142__A1 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09346__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17915_ net1603 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
X_13038_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[48\] net1933 net868 vssd1 vssd1
+ vccd1 vccd1 _02087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11982__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1150 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[17\] vssd1 vssd1 vccd1 vccd1
+ net1150 sky130_fd_sc_hd__buf_2
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13763__A net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1161 team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 net1161
+ sky130_fd_sc_hd__clkbuf_4
X_17846_ clknet_leaf_64_wb_clk_i _03522_ _01786_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[116\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout1172 net1173 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__buf_2
XANTENNA__08857__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1183 net1185 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__buf_4
Xfanout1194 net1204 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17060__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14989_ net1212 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__inv_2
X_17777_ clknet_leaf_78_wb_clk_i _03453_ _01717_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11283__A _07188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17993__1493 vssd1 vssd1 vccd1 vccd1 _17993__1493/HI net1493 sky130_fd_sc_hd__conb_1
X_16728_ clknet_leaf_28_wb_clk_i _02415_ _00711_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16659_ clknet_leaf_129_wb_clk_i _02346_ _00642_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08872__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09200_ net1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[17\] net889
+ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_1346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11208__A1 _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12956__A1 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09131_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[14\] net932 vssd1
+ vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12318__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08624__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10627__A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09062_ net1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[12\] net898
+ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__and3_1
XANTENNA__10431__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08013_ net1412 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold600 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold611 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[73\] vssd1 vssd1 vccd1 vccd1
+ net2227 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_25_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout206_A _07855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold622 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[8\] vssd1 vssd1 vccd1 vccd1 net2238
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold633 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold644 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[22\] vssd1 vssd1 vccd1 vccd1
+ net2260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11392__B1 _04466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold666 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold677 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12053__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09964_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[3\] net816 net803 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[3\]
+ _06299_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__a221o_1
Xhold699 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1115_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16158__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13133__A1 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[2\] net652 _05227_ _05244_
+ _05247_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__a2111o_1
XANTENNA__17403__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12988__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09895_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[5\] net820 net758 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__a22o_1
Xhold1300 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2916 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14769__A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13095__D net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1311 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2938 sky130_fd_sc_hd__dlygate4sd3_1
X_08846_ _05160_ _05183_ _05184_ _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__or4_1
XFILLER_0_97_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1333 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1344 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1355 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[31\] vssd1 vssd1 vccd1 vccd1
+ net2982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1377 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08777_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[0\] net901 vssd1
+ vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1388 team_01_WB.instance_to_wrap.cpu.f0.state\[8\] vssd1 vssd1 vccd1 vccd1 net3004
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1399 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[23\] vssd1 vssd1 vccd1 vccd1
+ net3015 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17553__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11447__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_135_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10655__C1 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09598__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ net550 _06398_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08933__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09329_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[24\] net692 net688 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[24\]
+ _05668_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12228__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08615__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14149__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12340_ net2218 net265 net428 vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08007__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12271_ net2879 net241 net435 vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14010_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[73\] _04235_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[113\]
+ _04294_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__a221o_1
X_11222_ net554 _06980_ _07132_ _07560_ _07561_ vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__o311ai_1
XANTENNA__13372__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10186__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09040__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__A _07696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ _06254_ _06255_ _06284_ _06409_ vssd1 vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_43_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09328__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[6\] net958 vssd1
+ vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__and3_1
XANTENNA__17083__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15961_ net1333 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__inv_2
X_11084_ _05729_ _06811_ _07344_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__or3b_1
XANTENNA__14679__A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13675__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10035_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[0\] net951 vssd1
+ vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__and3_1
X_14912_ net1241 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
X_17700_ clknet_leaf_101_wb_clk_i _03384_ _01641_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11686__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15892_ net1388 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__inv_2
XANTENNA__08677__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17631_ clknet_leaf_114_wb_clk_i _03316_ _01572_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14843_ net1197 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17562_ clknet_leaf_60_wb_clk_i _03249_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14774_ net1247 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11986_ net2559 net296 net474 vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16513_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[11\]
+ _00496_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13725_ _04109_ _04131_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[14\]
+ sky130_fd_sc_hd__nor2_1
X_10937_ _07067_ _07157_ net515 vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17493_ clknet_leaf_126_wb_clk_i _03180_ _01476_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09004__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12927__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16444_ clknet_leaf_8_wb_clk_i _02198_ _00427_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13656_ _03872_ _03876_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10868_ _06740_ _07112_ _06715_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_136_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_72_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12607_ net2980 net257 net396 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__mux2_1
XANTENNA__11550__B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16375_ clknet_leaf_67_wb_clk_i _02129_ _00358_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12138__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08606__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13587_ _03902_ _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10799_ _07137_ _07138_ net517 vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18114_ net1593 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
X_15326_ net1275 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__inv_2
X_12538_ net2102 net265 net403 vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11977__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18045_ net1545 vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__buf_2
XFILLER_0_124_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15257_ net1258 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12469_ net3032 net239 net411 vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14208_ net2317 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__17426__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09674__C net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15188_ net1267 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__inv_2
XANTENNA__09031__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14139_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[95\] _04240_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[127\]
+ _04423_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout409 _03564_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_39_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16450__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13493__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08700_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] net702 _05036_ _05039_
+ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_20_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12601__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09680_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[22\] net794 _06010_ _06012_
+ _06013_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_98_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08587__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08542__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_143_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_143_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08631_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 net597 vssd1 vssd1 vccd1 vccd1
+ _04971_ sky130_fd_sc_hd__nand2_1
X_17829_ clknet_leaf_71_wb_clk_i _03505_ _01769_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08562_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[19\] net919
+ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_102_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14091__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10637__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08493_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[23\] net677 _04809_
+ _04824_ _04769_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08845__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08753__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12048__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09114_ _05418_ _05453_ net602 vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_21_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10404__A2 _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11887__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09045_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[12\] net921
+ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1232_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09558__B1 _05897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08261__S net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold430 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[30\] vssd1 vssd1 vccd1 vccd1
+ net2057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[57\] vssd1 vssd1 vccd1 vccd1
+ net2068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout692_A _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold463 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] vssd1 vssd1 vccd1 vccd1
+ net2079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold485 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_117_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold496 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10523__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout910 net912 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout921 _04770_ vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout932 net933 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__buf_4
X_09947_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[3\] net968 vssd1
+ vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__and3_1
Xfanout943 net944 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13657__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout954 net956 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__buf_6
XANTENNA_fanout957_A _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 _04645_ vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12511__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout976 net977 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__clkbuf_4
X_09878_ _06217_ _06216_ vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_77_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout987 _04491_ vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1
+ net2746 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout998 net999 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__buf_1
XFILLER_0_137_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2757 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08928__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08829_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[1\] net903 vssd1
+ vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__and3_1
Xhold1152 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1163 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2779 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1174 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2790 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1185 _04128_ vssd1 vssd1 vccd1 vccd1 net2801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2812 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ net2743 net237 net487 vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14082__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13850__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11771_ net1889 net240 net495 vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__mux2_1
XANTENNA__08836__A2 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13847__A_N net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13290__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18063__1563 vssd1 vssd1 vccd1 vccd1 _18063__1563/HI net1563 sky130_fd_sc_hd__conb_1
XFILLER_0_90_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13510_ _03844_ _03948_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10722_ net534 _07010_ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__or2_2
X_14490_ net1387 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13441_ _05456_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 _03902_ sky130_fd_sc_hd__and2b_1
X_10653_ _04706_ net543 net537 _06992_ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10267__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12871__A_N net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16160_ clknet_leaf_98_wb_clk_i _01923_ _00148_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13372_ net1655 net830 _03838_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1
+ vccd1 vccd1 _01875_ sky130_fd_sc_hd__a22o_1
X_10584_ _06901_ _06917_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__or2_2
XFILLER_0_24_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09261__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15111_ net1300 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__inv_2
XANTENNA__11797__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12323_ net2777 net292 net432 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__mux2_1
XANTENNA__13578__A _03914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16091_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[13\]
+ _00079_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[13\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09549__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15042_ net1313 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__inv_2
X_12254_ net2121 net305 net441 vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__mux2_1
X_17992__1492 vssd1 vssd1 vccd1 vccd1 _17992__1492/HI net1492 sky130_fd_sc_hd__conb_1
XFILLER_0_43_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10714__B _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11205_ net374 net334 net333 vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__a21o_1
X_12185_ net2863 net311 net449 vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08772__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09791__A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11136_ _07469_ _07470_ _07475_ vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__a21bo_2
XANTENNA__08772__B2 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16993_ clknet_leaf_42_wb_clk_i _02680_ _00976_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15944_ net1335 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__inv_2
XANTENNA__12421__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10730__A _05115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ _07368_ _07405_ _04947_ net375 vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_34_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14202__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10018_ _06346_ _06349_ _06354_ _06357_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_30_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15875_ net1353 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10331__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14826_ net1276 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__inv_2
X_17614_ clknet_leaf_110_wb_clk_i _03299_ _01555_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14073__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14757_ net1219 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__inv_2
X_17545_ clknet_leaf_14_wb_clk_i _03232_ _01528_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13281__B1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11969_ net2165 net203 net471 vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13708_ team_01_WB.instance_to_wrap.cpu.c0.count\[1\] team_01_WB.instance_to_wrap.cpu.c0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__or2_1
X_17476_ clknet_leaf_52_wb_clk_i _03163_ _01459_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14688_ net1360 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09669__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08573__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16427_ clknet_leaf_109_wb_clk_i _02181_ _00410_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13639_ net727 _07308_ net983 vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16358_ clknet_leaf_69_wb_clk_i _02112_ _00341_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10398__A1 _06737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09252__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15309_ net1210 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_93_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16289_ clknet_leaf_61_wb_clk_i _02043_ _00272_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[12\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_93_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16816__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_11__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18028_ net1528 vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__buf_2
XFILLER_0_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout206 _07855_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_2
X_09801_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[14\] net800 _06139_
+ _06140_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout217 _07835_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_1
XANTENNA__10343__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09960__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout228 _07900_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_1
XANTENNA__16966__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07993_ net1119 vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__clkinv_4
Xfanout239 _07870_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_108_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13639__A2 _07308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09732_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[20\] net976
+ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__and3_1
XANTENNA__10640__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12331__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08748__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09206__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[22\] net973
+ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__and3_1
XANTENNA__08110__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout273_A _07866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[11\] net691 net674 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__a22o_1
X_09594_ net512 _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14064__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08279__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08545_ net1141 net619 net593 vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout440_A _07962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1182_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11822__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16346__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[23\] net878 vssd1
+ vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__and3_1
XANTENNA__09491__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout705_A _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14782__A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xwire618 _05331_ vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13575__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09243__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08987__D1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13398__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12506__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09028_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[9\] net680 _05340_ _05350_
+ _05361_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold260 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[121\] vssd1 vssd1 vccd1 vccd1
+ net1876 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10026__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold271 net132 vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold282 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold293 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[2\] vssd1 vssd1 vccd1 vccd1
+ net1909 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout740 net742 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout751 _04680_ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__buf_4
Xfanout762 _04674_ vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__buf_6
XFILLER_0_102_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12241__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13990_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[112\] _04255_ _04260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[56\]
+ _04272_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__a221o_1
Xfanout773 net774 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_8
Xfanout784 _04661_ vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__buf_4
Xfanout795 net797 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__buf_4
X_12941_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[10\] net1035 vssd1 vssd1 vccd1
+ vccd1 _03704_ sky130_fd_sc_hd__or2_1
XANTENNA__11365__B team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08020__A team_01_WB.instance_to_wrap.cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15660_ net1209 vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12872_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[31\] _03654_ net1030 vssd1
+ vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__mux2_1
X_14611_ net1348 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11823_ net1891 net293 net493 vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__mux2_1
X_15591_ net1328 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
XANTENNA__10696__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13263__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17330_ clknet_leaf_131_wb_clk_i _03017_ _01313_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14542_ net1335 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__inv_2
XANTENNA__08166__S net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11754_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[0\] _07438_ net718 vssd1 vssd1
+ vccd1 vccd1 _07940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_7__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ clknet_leaf_2_wb_clk_i _02948_ _01244_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10705_ _05805_ _05867_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14473_ net1373 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11685_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[14\] net717 vssd1 vssd1 vccd1
+ vccd1 _07885_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16212_ clknet_leaf_62_wb_clk_i net1628 _00200_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13566__A1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13424_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] _04949_ _03884_ vssd1
+ vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__nor3_1
XANTENNA__09786__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10636_ net336 _06919_ _06975_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__mux2_1
X_17192_ clknet_leaf_24_wb_clk_i _02879_ _01175_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09234__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16143_ clknet_leaf_98_wb_clk_i _01906_ _00131_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13355_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] net1064 team_01_WB.instance_to_wrap.cpu.f0.i\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12416__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10567_ net512 net511 net543 vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11320__S _07655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13101__A net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12306_ net2177 net267 net431 vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__mux2_1
X_16074_ clknet_leaf_119_wb_clk_i _01867_ _00062_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_0_51_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16989__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13286_ _03773_ _03771_ net828 net2869 vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_126_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10498_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[31\] net943
+ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__and3_1
X_15025_ net1291 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_127_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12237_ net2565 net271 net441 vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10001__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12168_ net2510 net245 net447 vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__mux2_1
XANTENNA__09952__C net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10552__A1 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16219__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11119_ net556 _07456_ _07458_ vssd1 vssd1 vccd1 vccd1 _07459_ sky130_fd_sc_hd__o21a_1
XANTENNA__12151__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12829__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12099_ net2294 net274 net457 vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__mux2_1
X_16976_ clknet_leaf_13_wb_clk_i _02663_ _00959_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15927_ net1409 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__inv_2
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_1
XANTENNA__14867__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11990__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ net1386 vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__inv_2
XANTENNA__14046__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08865__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12057__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14809_ net1304 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15789_ net1317 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08330_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[30\] net951 vssd1
+ vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__and3_1
X_17528_ clknet_leaf_25_wb_clk_i _03215_ _01511_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15698__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[20\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[12\]
+ net1038 vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17459_ clknet_leaf_137_wb_clk_i _03146_ _01442_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10338__C net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08192_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[89\] net1629 net1050 vssd1 vssd1
+ vccd1 vccd1 _03495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09225__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12326__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10240__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10791__B2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10073__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18062__1562 vssd1 vssd1 vccd1 vccd1 _18062__1562/HI net1562 sky130_fd_sc_hd__conb_1
XFILLER_0_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1028_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09933__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout488_A _07947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12061__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__A net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 _04474_
+ sky130_fd_sc_hd__inv_2
XANTENNA__08478__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09715_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[21\] net746 _06041_ _06042_
+ _06048_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout655_A _04817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1397_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[23\] net731 _05969_ _05973_
+ _05975_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_65_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10846__A2 _06921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14037__A2 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09577_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[25\] net813 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout822_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17991__1491 vssd1 vssd1 vccd1 vccd1 _17991__1491/HI net1491 sky130_fd_sc_hd__conb_1
XFILLER_0_93_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08528_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[18\] net915
+ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08459_ net1107 net1110 net1113 net1114 vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_107_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09102__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13548__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11470_ net367 _07762_ net2755 net875 vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09216__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08941__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10421_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[27\] net970
+ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__and3b_1
XFILLER_0_33_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12236__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10231__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13140_ net100 net850 net633 net2476 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__a22o_1
XANTENNA__12771__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10352_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[17\] net735 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__a22o_1
XANTENNA__08015__A _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13071_ net3113 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[23\] net861 vssd1 vssd1
+ vccd1 vccd1 _02054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10283_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[19\] net775 net760 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__a22o_1
X_12022_ net3089 net319 net470 vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__mux2_1
XANTENNA_input49_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16830_ clknet_leaf_45_wb_clk_i _02517_ _00813_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout570 _04520_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17637__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13973_ _04217_ _04222_ _04239_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__and3_4
X_16761_ clknet_leaf_58_wb_clk_i _02448_ _00744_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15712_ net1241 vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__inv_2
X_12924_ _04944_ net580 net362 vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__a21oi_2
X_16692_ clknet_leaf_12_wb_clk_i _02379_ _00675_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08685__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14028__A2 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12919__B net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12855_ net2321 net253 net379 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
X_15643_ net1179 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11806_ net1951 net267 net491 vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__mux2_1
X_15574_ net1198 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12786_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[14\] _07188_ net1027 vssd1 vssd1
+ vccd1 vccd1 _03619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09455__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17313_ clknet_leaf_41_wb_clk_i _03000_ _01296_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14525_ net1405 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11737_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[4\] net718 vssd1 vssd1 vccd1
+ vccd1 _07927_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09012__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17244_ clknet_leaf_32_wb_clk_i _02931_ _01227_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14456_ net1361 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11668_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] _07812_ vssd1 vssd1
+ vccd1 vccd1 _07872_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09947__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08851__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13407_ _03866_ _03867_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_3_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10619_ _06945_ _06958_ net529 vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__mux2_1
X_17175_ clknet_leaf_136_wb_clk_i _02862_ _01158_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12146__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire960 net961 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_2
X_14387_ net1305 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11599_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _07814_ vssd1 vssd1
+ vccd1 vccd1 _07816_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10222__B1 _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16126_ clknet_leaf_91_wb_clk_i _00007_ _00114_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_109_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12762__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13338_ _07682_ _03812_ _03813_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_1340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11985__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16057_ clknet_leaf_91_wb_clk_i _01850_ _00045_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_13269_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] net1062 _03754_ _03755_ net565
+ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__o311a_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15008_ net1241 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11722__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11286__A _07019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10190__A _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16191__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16959_ clknet_leaf_8_wb_clk_i _02646_ _00942_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_09500_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[29\] net944 vssd1
+ vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09431_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[28\] net692 net688 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[28\]
+ _05770_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09362_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[25\] net697 net656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[25\]
+ _05701_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08313_ net1146 net1148 net1151 net1153 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__and4b_2
XFILLER_0_117_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09293_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[22\] net915 vssd1
+ vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__and3_1
XANTENNA_11 _06589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _07858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08244_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[37\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[29\]
+ net1040 vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__mux2_1
XANTENNA_33 _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_44 _07900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_55 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_66 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12202__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ net2328 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[98\] net1043 vssd1 vssd1
+ vccd1 vccd1 _03512_ sky130_fd_sc_hd__mux2_1
XANTENNA__12056__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout403_A _03565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10365__A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1145_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10213__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12753__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10764__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11895__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1312_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09906__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
XANTENNA__16534__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput173 net173 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput184 net184 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XANTENNA__10516__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10970_ _06255_ _06410_ _07291_ _07309_ net344 vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__a311o_1
XANTENNA__09685__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08936__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ net1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[23\] net957
+ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12640_ net2132 net255 net392 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09437__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12571_ net2697 net263 net399 vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14310_ net1350 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11522_ net1711 net1158 net588 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1
+ vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15290_ net1189 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08671__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14241_ net1331 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__inv_2
XANTENNA__16064__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11453_ net1161 _04621_ _07669_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1
+ vccd1 vccd1 _07751_ sky130_fd_sc_hd__a31o_1
XANTENNA__10275__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire278 _07579_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_2
X_10404_ _06598_ _06604_ _06743_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__a21o_1
X_14172_ net1412 _04446_ _04447_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__nor3_1
X_11384_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] _07712_ vssd1 vssd1 vccd1 vccd1
+ _07713_ sky130_fd_sc_hd__nand2_1
X_13123_ net87 net846 net635 net1621 vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10335_ _06673_ _06674_ _06672_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13054_ net2564 net2376 net860 vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__mux2_1
X_17931_ net1433 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
X_10266_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[19\] net959
+ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1310 net1311 vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__clkbuf_4
X_12005_ net2223 net239 net467 vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__mux2_1
Xfanout1321 net1322 vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__buf_4
Xfanout1332 net1334 vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__buf_4
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17862_ clknet_leaf_82_wb_clk_i _03537_ _01802_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10197_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[8\] net959 vssd1
+ vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__and3_1
Xfanout1343 net1345 vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__buf_4
XANTENNA__11180__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1354 net1358 vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__buf_4
Xfanout1365 net1366 vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__buf_4
X_16813_ clknet_leaf_139_wb_clk_i _02500_ _00796_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1376 net1378 vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__buf_4
XANTENNA__09007__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1387 net1389 vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__buf_4
X_17793_ clknet_leaf_77_wb_clk_i net3150 _01733_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1398 net1399 vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_21_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15306__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16744_ clknet_leaf_23_wb_clk_i _02431_ _00727_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13956_ _04223_ _04231_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__nand2_4
XANTENNA__14210__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09676__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13209__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12907_ _05615_ net577 net361 vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__o21ba_1
X_13887_ _04193_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__inv_2
X_16675_ clknet_leaf_23_wb_clk_i _02362_ _00658_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15626_ net1276 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__inv_2
X_12838_ net3054 net214 net380 vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09428__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18061__1561 vssd1 vssd1 vccd1 vccd1 _18061__1561/HI net1561 sky130_fd_sc_hd__conb_1
XFILLER_0_51_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16407__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15557_ net1210 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__inv_2
X_12769_ net1621 net639 net609 _03607_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14508_ net1392 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__inv_2
X_15488_ net1243 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__inv_2
XANTENNA__08581__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
X_17227_ clknet_leaf_4_wb_clk_i _02914_ _01210_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
X_14439_ net1376 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput53 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput64 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
Xhold804 _03513_ vssd1 vssd1 vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
X_17158_ clknet_leaf_40_wb_clk_i _02845_ _01141_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold815 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold826 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09600__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17802__CLK clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10746__B2 _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold837 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16109_ clknet_leaf_91_wb_clk_i _01884_ _00097_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_17089_ clknet_leaf_42_wb_clk_i _02776_ _01072_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_09980_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[2\] _04634_ net774 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[2\]
+ _06319_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__a221o_1
XANTENNA__12604__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold859 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990__1490 vssd1 vssd1 vccd1 vccd1 _17990__1490/HI net1490 sky130_fd_sc_hd__conb_1
X_08931_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[6\] net911 vssd1
+ vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09364__B2 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08862_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[3\] net894 vssd1
+ vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1504 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net3120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1515 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1526 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08793_ _05120_ _05124_ _05128_ _05132_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__or4_1
Xhold1537 team_01_WB.instance_to_wrap.a1.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net3153
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1548 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1559 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3175 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09116__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08756__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout353_A _03741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1095_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[27\] net693 net676 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[27\]
+ _05740_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__a221o_1
XANTENNA__10682__A0 _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[25\] net937
+ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout520_A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10434__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09276_ net1116 net713 net594 vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08227_ net2394 net2668 net1038 vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09884__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08158_ net1643 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[115\] net1052 vssd1 vssd1
+ vccd1 vccd1 _03529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17482__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout987_A _04491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08089_ _04523_ _04530_ _04536_ _04542_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__or4_2
XFILLER_0_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12514__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10120_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[6\] net787 _04667_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[6\]
+ _06459_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11638__B _07600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10051_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[0\] net802 net790 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13853__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11654__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ net3095 net833 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[3\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_19_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14790_ net1292 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09124__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13741_ net1165 net1855 net1054 vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__a21o_1
X_10953_ _06441_ _06470_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16460_ clknet_leaf_142_wb_clk_i _02214_ _00443_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13672_ net1649 net567 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1
+ vccd1 vccd1 _01830_ sky130_fd_sc_hd__a22o_1
X_10884_ net335 _07222_ _07223_ net337 vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08963__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15411_ net1280 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12623_ net2365 net225 net391 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__mux2_1
X_16391_ clknet_leaf_67_wb_clk_i net2726 _00374_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08618__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15342_ net1282 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__inv_2
XANTENNA__10425__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12965__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12554_ net2813 net291 net404 vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__mux2_1
XANTENNA__08174__S net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10976__A1 _07015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09830__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[10\] _07756_ vssd1 vssd1 vccd1
+ vccd1 _07780_ sky130_fd_sc_hd__and2_1
X_15273_ net1230 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__inv_2
X_18061_ net1561 vssd1 vssd1 vccd1 vccd1 la_data_out[103] sky130_fd_sc_hd__buf_2
X_12485_ net2231 net305 net414 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14224_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] vssd1 vssd1 vccd1
+ vccd1 _02263_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09794__A _06129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17012_ clknet_leaf_13_wb_clk_i _02699_ _00995_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11436_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] _07736_ _07742_ vssd1 vssd1 vccd1
+ vccd1 _03372_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12932__B net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14155_ net1782 _04195_ net1411 vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12424__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367_ _04575_ _07651_ vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__or2_2
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13106_ net637 vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__inv_2
X_10318_ net987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[18\] net941 vssd1
+ vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__o21a_1
X_14086_ _04367_ _04369_ _04371_ _04373_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11548__B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11298_ net1068 _07637_ vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13037_ net2786 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[57\] net866 vssd1 vssd1
+ vccd1 vccd1 _02088_ sky130_fd_sc_hd__mux2_1
XANTENNA__13142__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17914_ net1430 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XFILLER_0_123_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10249_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[9\] net766 _06583_ _06588_
+ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__o22a_2
XFILLER_0_119_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09897__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1140 net1141 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__clkbuf_2
Xfanout1151 net1152 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__clkbuf_2
X_17845_ clknet_leaf_73_wb_clk_i _03521_ _01785_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[115\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1162 team_01_WB.instance_to_wrap.cpu.f0.state\[4\] vssd1 vssd1 vccd1 vccd1
+ net1162 sky130_fd_sc_hd__buf_2
Xfanout1173 net1204 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__buf_4
Xfanout1184 net1185 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__buf_4
XANTENNA__15036__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1195 net1203 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__buf_4
X_17776_ clknet_leaf_86_wb_clk_i net2669 _01716_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_14988_ net1206 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__inv_2
XANTENNA__09649__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16727_ clknet_leaf_138_wb_clk_i _02414_ _00710_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11283__B _07232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13939_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__nor2_2
XFILLER_0_92_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12653__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16658_ clknet_leaf_129_wb_clk_i _02345_ _00641_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15609_ net1260 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08609__B1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16589_ clknet_leaf_138_wb_clk_i _02276_ _00572_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13602__B1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09130_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[14\] net914 vssd1
+ vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10967__A1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10627__B net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09061_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[12\] net912
+ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_117_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09200__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08012_ net1 vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__inv_2
XANTENNA__10346__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire955_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold601 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold612 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold623 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold634 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12334__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold645 team_01_WB.instance_to_wrap.a1.ADR_I\[14\] vssd1 vssd1 vccd1 vccd1 net2261
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11392__A1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_107_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09963_ _06286_ _06300_ _06301_ _06302_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__or4_1
XANTENNA__13669__A0 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11458__B net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold678 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09209__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold689 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_65_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08914_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[2\] net659 _05243_ _05245_
+ net708 vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13133__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[5\] net801 net783 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1010_A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1301 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[65\] vssd1 vssd1 vccd1 vccd1
+ net2917 sky130_fd_sc_hd__dlygate4sd3_1
X_08845_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[1\] net663 net658 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__a22o_1
Xhold1312 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1323 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1334 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1345 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1356 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1367 _02070_ vssd1 vssd1 vccd1 vccd1 net2983 sky130_fd_sc_hd__dlygate4sd3_1
X_08776_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] _04751_ _04752_ net1116 vssd1
+ vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__a22o_2
XANTENNA__14094__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1378 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1389 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3005 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08486__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11193__B net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout735_A _04687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout902_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12509__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09328_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[24\] net701 net656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold313_A team_01_WB.instance_to_wrap.cpu.f0.write_data\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09273__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09812__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10958__A1 _05042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11080__B1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09259_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[20\] net681 net677 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[20\]
+ _05596_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16872__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09818__S net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12270_ net3249 net273 net437 vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__mux2_1
XANTENNA__13848__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ net554 _07202_ _07017_ vssd1 vssd1 vccd1 vccd1 _07561_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11649__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13372__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12244__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__A2 _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09119__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _06284_ _06409_ _06254_ _06255_ vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__o211a_1
XANTENNA__17228__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10103_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[6\] net979 vssd1
+ vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__and3_1
X_15960_ net1336 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__inv_2
X_11083_ _05681_ net511 _07349_ _05707_ net512 vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__o32a_1
XFILLER_0_60_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18060__1560 vssd1 vssd1 vccd1 vccd1 _18060__1560/HI net1560 sky130_fd_sc_hd__conb_1
XANTENNA__11135__B2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[0\] net948 vssd1
+ vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__and3_1
X_14911_ net1257 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15891_ net1397 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__inv_2
XANTENNA__12883__A1 _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11686__A2 _07188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11384__A team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17630_ clknet_leaf_118_wb_clk_i _03315_ _01571_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_51_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ net1190 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14085__B1 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08169__S net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17561_ clknet_leaf_60_wb_clk_i _03248_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11985_ net2807 net301 net474 vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__mux2_1
X_14773_ net1219 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10646__A0 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16512_ clknet_leaf_112_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[10\]
+ _00495_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10936_ net556 _07069_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13724_ net3288 _04108_ net1972 vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__a21oi_1
X_17492_ clknet_leaf_128_wb_clk_i _03179_ _01475_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10110__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16443_ clknet_leaf_46_wb_clk_i _02197_ _00426_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10867_ _07205_ _07206_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__or2_2
XANTENNA__12419__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13655_ net983 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] _04087_ _04088_
+ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10728__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12606_ net2073 net260 net396 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__mux2_1
X_16374_ clknet_leaf_69_wb_clk_i _02128_ _00357_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09264__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13586_ _03912_ _04029_ _03903_ _03906_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10798_ net513 _05898_ net504 _06811_ net548 net538 vssd1 vssd1 vccd1 vccd1 _07138_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09803__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18113_ net638 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15325_ net1253 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__inv_2
X_12537_ net1999 net268 net403 vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__mux2_1
XANTENNA__09020__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18044_ net1544 vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__buf_2
X_12468_ net3138 net272 net413 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__mux2_1
X_15256_ net1178 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09955__C net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11419_ _04478_ _07702_ vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__nand2_1
X_14207_ net2809 vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__clkbuf_1
X_15187_ net1281 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__inv_2
XANTENNA__12154__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12399_ net2953 net208 net419 vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14138_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[127\] _04263_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11993__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14069_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[92\] _04240_ _04249_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__a22o_1
XANTENNA__12874__A1 _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08542__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08630_ net377 vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__inv_2
X_17828_ clknet_leaf_66_wb_clk_i _03504_ _01768_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14076__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08561_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[19\] net934
+ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__and3_1
X_17759_ clknet_leaf_64_wb_clk_i _03435_ _01699_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[29\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_76_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09699__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08492_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[23\] net697 _04802_
+ _04805_ _04814_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_112_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12329__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08108__A _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09113_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] net703 _05449_ _05452_
+ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout316_A _07939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1058_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10076__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[12\] net933
+ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__and3_1
XANTENNA__16125__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14000__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09558__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold420 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[16\] vssd1 vssd1 vccd1 vccd1 net2036
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12064__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold431 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[5\] vssd1 vssd1 vccd1 vccd1
+ net2047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10168__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold442 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1225_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold453 _03471_ vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold464 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 net2080
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[59\] vssd1 vssd1 vccd1 vccd1
+ net2091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold486 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16275__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout685_A _04780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout900 net905 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold497 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 net912 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__buf_4
Xfanout922 net924 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09946_ net993 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[3\] net955 vssd1
+ vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_70_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout933 _04762_ vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_8
XANTENNA__17520__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout944 _04665_ vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13511__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout966 net968 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__buf_4
XFILLER_0_99_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1120 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[96\] vssd1 vssd1 vccd1 vccd1
+ net2736 sky130_fd_sc_hd__dlygate4sd3_1
X_09877_ _05416_ _06189_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_5_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout988 net990 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__buf_2
Xhold1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2747 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08533__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout999 net1014 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__buf_2
Xhold1142 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[11\] vssd1 vssd1 vccd1 vccd1
+ net2758 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ net1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[1\] net890 vssd1
+ vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__and3_1
Xhold1153 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2769 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2780 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1175 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2791 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2802 sky130_fd_sc_hd__dlygate4sd3_1
X_08759_ net1088 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[4\] net923 vssd1
+ vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1197 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2813 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17670__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10628__A0 _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11770_ net2463 _07866_ net497 vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10721_ _07006_ _07013_ net534 vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__mux2_1
XANTENNA__08944__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12239__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11143__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13440_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _04945_ vssd1 vssd1
+ vccd1 vccd1 _03901_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10652_ net548 net513 vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09246__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13371_ net585 net564 net826 vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_131_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10583_ _06901_ _06917_ vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12322_ net3156 net316 net434 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__mux2_1
X_15110_ net1293 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16090_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[12\]
+ _00078_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[12\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17050__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15041_ net1246 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__inv_2
X_12253_ net2293 net309 net440 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__mux2_1
X_11204_ _06218_ _07173_ _06194_ vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12184_ net2090 net295 net449 vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11135_ _07040_ _07338_ _07471_ net345 _07474_ vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_53_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12702__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16992_ clknet_leaf_32_wb_clk_i _02679_ _00975_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15943_ net1409 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__inv_2
X_11066_ _05491_ _06158_ _07366_ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_34_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10017_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[1\] net759 _06355_ _06356_
+ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14058__B1 _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15874_ net1330 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17613_ clknet_leaf_79_wb_clk_i _03298_ _01554_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14825_ net1229 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__inv_2
XANTENNA__09015__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15314__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17544_ clknet_leaf_22_wb_clk_i _03231_ _01527_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09485__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14756_ net1345 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__inv_2
XANTENNA__13281__A1 _07650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ net1808 net205 net471 vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08854__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13707_ net1994 _04100_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[2\]
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_47_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10919_ _05374_ net340 vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__xnor2_2
X_17475_ clknet_leaf_20_wb_clk_i _03162_ _01458_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12149__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11899_ net2723 net210 net481 vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__mux2_1
X_14687_ net1365 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13569__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16426_ clknet_leaf_106_wb_clk_i _02180_ _00409_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16148__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09237__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13638_ net188 _04073_ _04074_ net727 vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11988__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16357_ clknet_leaf_74_wb_clk_i _02111_ _00340_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13569_ net186 _04015_ _04016_ net726 vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15308_ net1197 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_93_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16288_ clknet_leaf_73_wb_clk_i _02042_ _00271_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16298__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18027_ net1527 vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__buf_2
XANTENNA__11289__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15239_ net1328 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09800_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[14\] _04667_ net735
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[14\] vssd1 vssd1 vccd1 vccd1
+ _06140_ sky130_fd_sc_hd__a22o_1
XANTENNA__08763__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout207 net208 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__buf_2
Xfanout218 _07835_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_2
X_07992_ net1084 vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__inv_2
XANTENNA__12612__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout229 _07900_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_2
XFILLER_0_5_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09731_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[20\] net970
+ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10640__B _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10858__A0 _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09662_ _05999_ _06000_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__nand2_1
XANTENNA__14049__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08613_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[11\] net682 net669 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__a22o_1
X_09593_ _05707_ _05735_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout266_A _07880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08544_ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__inv_2
XANTENNA__09476__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11471__B net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08475_ net1007 net879 vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__and2_1
XANTENNA__12059__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout433_A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10368__A _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1175_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_59_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11898__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout600_A _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1342_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10389__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08272__S net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_80_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09027_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[9\] _04771_ _05344_ _05353_
+ _05355_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__a2111o_1
XANTENNA__15894__A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09892__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold250 _02016_ vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 _03527_ vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold272 _01997_ vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 net112 vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold294 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout741 net742 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__buf_6
XANTENNA__08939__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09929_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[4\] net821 net790 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__a22o_1
Xfanout752 _04678_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__buf_6
Xfanout763 _04674_ vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout774 _04669_ vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_8
Xfanout785 net786 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__buf_6
Xfanout796 net797 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_6
X_12940_ net584 _07757_ _03694_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12871_ net873 team_01_WB.instance_to_wrap.cpu.RU0.next_write_i vssd1 vssd1 vccd1
+ vccd1 _03655_ sky130_fd_sc_hd__and2b_1
X_14610_ net1348 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__inv_2
X_11822_ net2332 net316 net494 vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__mux2_1
X_15590_ net1299 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
XANTENNA__13263__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09467__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09132__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08674__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11753_ net2773 net316 net502 vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__mux2_1
X_14541_ net1394 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10278__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09482__A3 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10704_ _05806_ net513 vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__nor2_1
X_17260_ clknet_leaf_133_wb_clk_i _02947_ _01243_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14472_ net1336 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11684_ net2405 net232 net500 vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16211_ clknet_leaf_62_wb_clk_i net1838 _00199_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13423_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] net1156 net730 _04838_ net1116
+ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__a32o_1
XANTENNA__13566__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10635_ _04707_ _05835_ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17191_ clknet_leaf_15_wb_clk_i _02878_ _01174_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17566__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16142_ clknet_leaf_96_wb_clk_i _01905_ _00130_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13354_ net1706 _03826_ net826 vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__mux2_1
XANTENNA__08182__S net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10566_ net525 net519 vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__nand2_4
XFILLER_0_84_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12305_ net2994 net235 net431 vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13285_ _04621_ _03753_ _03772_ net828 vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__o31a_1
X_16073_ clknet_leaf_120_wb_clk_i _01866_ _00061_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\]
+ sky130_fd_sc_hd__dfstp_2
X_10497_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[31\] net799 net782 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10444__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11329__B2 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15024_ net1226 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__inv_2
X_12236_ net3273 net243 net439 vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16590__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15309__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12432__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ net2011 net203 net447 vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__mux2_1
XANTENNA__14213__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11118_ _06928_ _07133_ _07457_ net330 vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__a211o_1
XANTENNA__12829__A1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16975_ clknet_leaf_141_wb_clk_i _02662_ _00958_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12098_ net2652 net209 net457 vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15926_ net1395 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__inv_2
X_11049_ net520 _06339_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_1
XANTENNA__10304__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15857_ net1367 vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14808_ net1178 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09458__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15788_ net1315 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__inv_2
XANTENNA__08584__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17527_ clknet_leaf_140_wb_clk_i _03214_ _01510_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14739_ net1308 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__inv_2
XANTENNA__10188__A _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[21\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[13\]
+ net1040 vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17458_ clknet_leaf_134_wb_clk_i _03145_ _01441_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_95_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08881__A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16409_ clknet_leaf_61_wb_clk_i _02163_ _00392_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08191_ net2245 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[82\] net1043 vssd1 vssd1
+ vccd1 vccd1 _03496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12607__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17389_ clknet_leaf_2_wb_clk_i _03076_ _01372_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11511__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16933__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10635__B _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08984__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08736__A2 _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13190__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15219__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12342__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08759__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 _04473_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout383_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09714_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[21\] net811 net772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[21\]
+ _06053_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09645_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[23\] net818 net791 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[23\]
+ _05984_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout550_A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1292_A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A _04825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09576_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[25\] net803 _05904_
+ _05911_ _05913_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09449__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13245__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08527_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[18\] net907
+ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout815_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16463__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09887__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[23\] net889
+ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13548__A2 _07154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12517__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08389_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\] _04623_ _04626_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_107_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10420_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[27\] net942
+ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12756__B1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08975__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10351_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[17\] net819 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_76_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13070_ net1783 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[24\] net860 vssd1 vssd1
+ vccd1 vccd1 _02055_ sky130_fd_sc_hd__mux2_1
X_10282_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[19\] net818 net772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12021_ net2182 net307 net470 vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08727__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12252__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__A _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10534__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08669__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout560 net561 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_2
Xfanout571 _04196_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14130__C1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16760_ clknet_leaf_27_wb_clk_i _02447_ _00743_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13972_ _04222_ _04237_ _04239_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__and3_4
Xfanout593 _04845_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08966__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15711_ net1260 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__inv_2
XANTENNA__10298__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ net2036 net871 net358 _03691_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16691_ clknet_leaf_135_wb_clk_i _02378_ _00674_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_85_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15642_ net1191 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12854_ net2677 net228 net381 vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11805_ net2557 net235 net491 vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15573_ net1222 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__inv_2
XANTENNA_output100_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12785_ net1771 net640 net607 _03618_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17312_ clknet_leaf_29_wb_clk_i _02999_ _01295_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14524_ net1392 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__inv_2
XANTENNA__09797__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11736_ net1827 net294 net501 vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16956__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12935__B net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17243_ clknet_leaf_17_wb_clk_i _02930_ _01226_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14455_ net1344 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12427__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[18\] _07251_ net716 vssd1 vssd1
+ vccd1 vccd1 _07871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13406_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] net595 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__a21o_1
X_10618_ _06950_ _06957_ net520 vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__mux2_1
X_17174_ clknet_leaf_141_wb_clk_i _02861_ _01157_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14386_ net1304 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11598_ _07814_ vssd1 vssd1 vccd1 vccd1 _07815_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10222__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16125_ clknet_leaf_5_wb_clk_i _00025_ _00113_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dfrtp_1
X_10549_ net510 net509 net543 vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__mux2_1
X_13337_ net1065 _07682_ _03811_ _04518_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__a211o_1
XFILLER_0_40_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16056_ clknet_leaf_92_wb_clk_i _01849_ _00044_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_122_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13268_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] _03749_ vssd1 vssd1 vccd1 vccd1
+ _03759_ sky130_fd_sc_hd__or2_1
XANTENNA__13172__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15007_ net1255 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12219_ net2831 net306 net445 vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__mux2_1
XANTENNA__12162__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13199_ net9 net835 net628 net2338 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_88_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11722__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11286__B _07056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08298__D net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16958_ clknet_leaf_46_wb_clk_i _02645_ _00941_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09143__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15909_ net1408 vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16889_ clknet_leaf_51_wb_clk_i _02576_ _00872_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_09430_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[28\] net700 net655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13227__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09361_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[25\] net672 net668 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[25\]
+ _05685_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__a221o_1
XANTENNA__09203__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08312_ net1131 net979 vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_19_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10349__C net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09292_ net1073 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[22\] net915
+ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_12 _06589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08243_ net3221 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[30\] net1037 vssd1 vssd1
+ vccd1 vccd1 _03444_ sky130_fd_sc_hd__mux2_1
XANTENNA__17881__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09500__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _07858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12337__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_45 _07900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A _07900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_56 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_67 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08174_ net2419 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[99\] net1052 vssd1 vssd1
+ vccd1 vccd1 _03513_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_127_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08116__A team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08957__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17111__CLK clknet_leaf_137_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1040_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10764__A2 _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1138_A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_88_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XANTENNA__13163__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput174 net174 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12072__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11713__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17261__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__A2 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08590__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16829__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout932_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09628_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[23\] net794 net740 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17939__1439 vssd1 vssd1 vccd1 vccd1 _17939__1439/HI net1439 sky130_fd_sc_hd__conb_1
XFILLER_0_112_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09559_ _05898_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12570_ net2035 net268 net399 vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09842__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16209__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11521_ net1158 _07784_ vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__nor2_1
XANTENNA__12247__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14240_ net1349 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__inv_2
X_11452_ _07672_ _07750_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10403_ _06641_ _06677_ _06715_ _06742_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__or4_1
X_14171_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[7\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\]
+ _04189_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__and3_1
XANTENNA__11401__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11383_ net1063 _07700_ _07710_ vssd1 vssd1 vccd1 vccd1 _07712_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13122_ net88 net844 net635 net1848 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a22o_1
X_10334_ net559 _05568_ _04883_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__o21ai_1
XANTENNA_input61_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13154__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13053_ net3176 net2922 net866 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11387__A _04466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17930_ net1432 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
X_10265_ net1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[19\] net941
+ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10291__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1300 net1301 vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__buf_4
XANTENNA__12901__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12004_ net2028 net273 net469 vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__mux2_1
Xfanout1311 net1314 vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__buf_4
X_17861_ clknet_leaf_82_wb_clk_i _03536_ _01801_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09373__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[8\] net949 vssd1
+ vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__and3_1
Xfanout1322 net1342 vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__buf_2
Xfanout1333 net1334 vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__buf_4
Xfanout1344 net1345 vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__buf_4
XFILLER_0_108_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16812_ clknet_leaf_133_wb_clk_i _02499_ _00795_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1355 net1358 vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__clkbuf_4
Xfanout1366 net1369 vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__buf_4
XANTENNA__12710__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17792_ clknet_leaf_65_wb_clk_i net2395 _01732_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_91_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1377 net1378 vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__buf_4
Xfanout1388 net1389 vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__clkbuf_4
Xfanout390 _03569_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_6
Xfanout1399 net1404 vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16743_ clknet_leaf_16_wb_clk_i _02430_ _00726_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13955_ _04219_ _04222_ _04237_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__and3_4
X_12906_ net2639 net871 net358 _03679_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__a22o_1
X_16674_ clknet_leaf_34_wb_clk_i _02361_ _00657_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13209__A1 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08884__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13886_ _04190_ _04191_ _04192_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__or3_2
XANTENNA__10140__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08884__B2 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15625_ net1229 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12837_ net2143 net217 net380 vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15556_ net1240 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__inv_2
XANTENNA__09833__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12768_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] net1055 net363 _03606_
+ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__a22o_1
XANTENNA__08862__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14507_ net1407 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11719_ net1949 net304 net501 vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15487_ net1257 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__inv_2
XANTENNA__17134__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12699_ net2785 _07866_ net385 vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17226_ clknet_leaf_11_wb_clk_i _02913_ _01209_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14438_ net1396 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__inv_2
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_1
XFILLER_0_71_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput43 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11996__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput54 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
X_17157_ clknet_leaf_32_wb_clk_i _02844_ _01140_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput65 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
X_14369_ net1343 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold805 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold816 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_137_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_137_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16108_ clknet_leaf_91_wb_clk_i _01883_ _00096_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold827 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17284__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold838 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[46\] vssd1 vssd1 vccd1 vccd1
+ net2465 sky130_fd_sc_hd__dlygate4sd3_1
X_17088_ clknet_leaf_29_wb_clk_i _02775_ _01071_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13145__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16039_ clknet_leaf_68_wb_clk_i _01833_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_08930_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[6\] net921 vssd1
+ vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08861_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[3\] net924 vssd1
+ vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__and3_1
Xhold1505 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1516 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08792_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[0\] net672 _05129_ _05130_
+ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12620__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1527 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1538 team_01_WB.instance_to_wrap.cpu.f0.num\[7\] vssd1 vssd1 vccd1 vccd1 net3154
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1549 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09413_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[27\] net678 net654 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[27\]
+ _05739_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__a221o_1
XANTENNA__10682__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout346_A net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10079__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12959__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[25\] net904
+ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13620__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09230__A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09275_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\] net704 _05610_ _05614_
+ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__o22a_2
XFILLER_0_69_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12067__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_136_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout513_A _05867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1255_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08226_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[55\] net2003 net1047 vssd1 vssd1
+ vccd1 vccd1 _03461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17627__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08157_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[124\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[116\]
+ net1041 vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08088_ _04525_ _04559_ _04560_ net569 team_01_WB.instance_to_wrap.cpu.f0.write_data\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__a32o_1
XFILLER_0_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout882_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13136__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17777__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10050_ _06386_ _06387_ _06388_ _06389_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__or4_1
XANTENNA__09355__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15407__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12530__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08947__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14100__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13740_ net1165 net1061 net1618 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__a21o_1
XANTENNA__10122__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ _06255_ _06410_ _07291_ _06468_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13671_ net1675 net567 net346 team_01_WB.instance_to_wrap.cpu.f0.i\[30\] vssd1 vssd1
+ vccd1 vccd1 _01831_ sky130_fd_sc_hd__a22o_1
XANTENNA__17157__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10883_ _05566_ _06707_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__xnor2_1
X_15410_ net1235 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__inv_2
XANTENNA__15142__A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12622_ net3216 net190 net391 vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__mux2_1
X_16390_ clknet_leaf_68_wb_clk_i net1746 _00373_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09815__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08682__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15341_ net1212 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12553_ net3009 net317 net406 vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10976__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18060_ net1560 vssd1 vssd1 vccd1 vccd1 la_data_out[102] sky130_fd_sc_hd__buf_2
X_11504_ net1635 net876 _07758_ _07779_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__o22a_1
X_15272_ net1288 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ net2387 net310 net412 vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17011_ clknet_leaf_135_wb_clk_i _02698_ _00994_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14223_ net3180 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11435_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] _07736_ net326 vssd1 vssd1 vccd1
+ vccd1 _07742_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12705__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14154_ net1714 net605 _04437_ net1170 vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__o211a_1
X_11366_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] team_01_WB.instance_to_wrap.cpu.f0.i\[23\]
+ net1063 _07694_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__and4_1
XANTENNA__10733__B _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13127__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10317_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[18\] net731 _06654_ _06655_
+ _06656_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__a2111o_1
X_13105_ _03723_ _03724_ _03725_ _03728_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__or4_1
X_14085_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[100\] _04254_ _04265_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\]
+ _04372_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__a221o_1
X_11297_ net199 net195 net615 vssd1 vssd1 vccd1 vccd1 _07637_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10452__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09346__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13036_ net2300 net2192 net857 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__mux2_1
X_10248_ net771 _06572_ _06575_ _06587_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__or4_1
X_17913_ net1429 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XFILLER_0_24_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09018__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1130 net1132 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_119_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1141 net1142 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__clkbuf_4
X_17844_ clknet_leaf_65_wb_clk_i _03520_ _01784_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_10179_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[10\] net795 net761 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[10\]
+ _06518_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__a221o_1
Xfanout1152 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1 vccd1
+ net1152 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12440__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1163 net1164 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__clkbuf_2
Xfanout1174 net1177 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__buf_4
Xfanout1185 net1204 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__buf_2
XANTENNA__08857__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17775_ clknet_leaf_62_wb_clk_i _03451_ _01715_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[45\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_89_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1196 net1203 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__buf_2
X_14987_ net1296 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__inv_2
X_16726_ clknet_leaf_141_wb_clk_i _02413_ _00709_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13938_ _04225_ _04229_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__nor2_8
XANTENNA__11283__C _07553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16657_ clknet_leaf_18_wb_clk_i _02344_ _00640_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13869_ net1164 net1059 net2078 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[30\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_69_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11580__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13271__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18009__1509 vssd1 vssd1 vccd1 vccd1 _18009__1509/HI net1509 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_100_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15608_ net1188 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09806__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16588_ clknet_leaf_117_wb_clk_i _02275_ _00571_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13602__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15539_ net1281 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__inv_2
XANTENNA__15987__A net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11613__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09060_ net1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[12\] net904
+ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08011_ team_01_WB.instance_to_wrap.a1.READ_I vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17209_ clknet_leaf_58_wb_clk_i _02896_ _01192_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09034__A1 _05373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16674__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12615__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold602 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[18\] vssd1 vssd1 vccd1 vccd1
+ net2229 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13300__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold624 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap343 _05378_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold635 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold646 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[70\] vssd1 vssd1 vccd1 vccd1
+ net2262 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13118__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold657 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
X_17938__1438 vssd1 vssd1 vccd1 vccd1 _17938__1438/HI net1438 sky130_fd_sc_hd__conb_1
Xhold668 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold679 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09962_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[3\] net801 net792 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08913_ _05249_ _05250_ _05251_ _05252_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__or4_1
XFILLER_0_110_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09893_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[5\] net950 vssd1
+ vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout296_A _07926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08545__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1302 _02096_ vssd1 vssd1 vccd1 vccd1 net2918 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12350__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[1\] net653 _05165_ _05169_
+ _05172_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__a2111o_1
Xhold1313 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2929 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10352__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1003_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1324 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1357 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2973 sky130_fd_sc_hd__dlygate4sd3_1
X_08775_ net599 _05110_ _05113_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_79_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1368 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2984 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout463_A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1379 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2995 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_0_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10655__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1372_A net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_40_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout728_A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09598__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09327_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[24\] net666 net663 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[24\]
+ _05666_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_62_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10958__A2 _06924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14149__A2 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11080__A1 _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09258_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[20\] net701 net670 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08209_ net2881 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[64\] net1049 vssd1 vssd1
+ vccd1 vccd1 _03478_ sky130_fd_sc_hd__mux2_1
XANTENNA__12525__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09189_ _05495_ _05528_ net600 vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__mux2_2
XFILLER_0_107_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ net369 _07343_ _07344_ net336 _07559_ vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__o221a_1
XFILLER_0_121_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09576__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08304__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ _07449_ net322 _07490_ vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10102_ _06441_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__inv_2
XANTENNA__09328__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11082_ _04844_ _05997_ _07418_ _07419_ _07421_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_120_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10033_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[0\] net815 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__a22o_1
X_14910_ net1248 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
XANTENNA__12260__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15890_ net1383 vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__inv_2
XANTENNA__09135__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08677__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ net1258 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ clknet_leaf_60_wb_clk_i _03247_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_14772_ net1267 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__inv_2
XANTENNA__08974__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11984_ net2043 net282 net471 vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16511_ clknet_leaf_112_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[9\]
+ _00494_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10646__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13723_ net2159 _04108_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[13\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_105_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10935_ net556 _07069_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17491_ clknet_leaf_136_wb_clk_i _03178_ _01474_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16442_ clknet_leaf_19_wb_clk_i _02196_ _00425_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08185__S net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13654_ net728 _07449_ net983 vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__a21oi_1
X_10866_ net563 _07192_ _07193_ _07203_ net558 vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13596__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12605_ net2679 net233 net397 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16373_ clknet_leaf_76_wb_clk_i _02127_ _00356_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13585_ _03912_ _04029_ _03906_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09301__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10797_ net512 net511 net510 net509 net548 net537 vssd1 vssd1 vccd1 vccd1 _07137_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_121_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10447__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18112_ net638 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15324_ net1174 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__inv_2
X_12536_ net2692 net235 net403 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18043_ net1543 vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__buf_2
XFILLER_0_87_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15255_ net1199 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__inv_2
X_12467_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[21\] net244 net411 vssd1
+ vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__mux2_1
XANTENNA__12435__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14206_ net3222 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__clkbuf_1
X_11418_ _07691_ _07732_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15186_ net1232 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__inv_2
X_12398_ net2769 net277 net422 vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14137_ _04416_ _04417_ _04419_ _04421_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_91_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11349_ team_01_WB.instance_to_wrap.cpu.f0.i\[11\] _07677_ vssd1 vssd1 vccd1 vccd1
+ _07678_ sky130_fd_sc_hd__nand2_2
X_14068_ net148 net605 vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__or2_1
XANTENNA__13870__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11575__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13019_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[67\] net1976 net865 vssd1 vssd1
+ vccd1 vccd1 _02106_ sky130_fd_sc_hd__mux2_1
XANTENNA__12170__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12874__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08587__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17827_ clknet_leaf_68_wb_clk_i _03503_ _01767_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14886__A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13790__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08560_ _04889_ _04893_ _04895_ _04899_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__or4_1
X_17758_ clknet_leaf_56_wb_clk_i _03434_ _01698_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[28\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_102_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17472__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10637__A1 _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16709_ clknet_leaf_38_wb_clk_i _02396_ _00692_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_08491_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[23\] net670 _04812_ _04820_
+ _04798_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17689_ clknet_leaf_99_wb_clk_i _03373_ _01630_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10919__A _05374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11514__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09255__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09211__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08108__B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09112_ _05443_ _05444_ _05450_ _05451_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_21_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09043_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[12\] net905
+ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14000__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12345__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout211_A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout309_A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold410 _02020_ vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09558__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11469__B net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold421 _01982_ vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold432 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold443 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12562__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold454 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1159_A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1120_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold465 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 _02098_ vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1218_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold487 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold498 team_01_WB.instance_to_wrap.cpu.f0.num\[22\] vssd1 vssd1 vccd1 vccd1 net2114
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout901 net902 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__clkbuf_4
X_09945_ _06280_ _06283_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__nand2_1
Xfanout912 _04779_ vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout923 net924 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_4
Xfanout934 net936 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout945 net947 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout678_A _04790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12080__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09876_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _06215_ net624 vssd1
+ vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__mux2_2
Xfanout967 net968 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__buf_2
Xhold1110 _02145_ vssd1 vssd1 vccd1 vccd1 net2726 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout978 net979 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_8
Xhold1121 _02135_ vssd1 vssd1 vccd1 vccd1 net2737 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 net990 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2748 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08827_ net1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[1\] net898 vssd1
+ vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__and3_1
XANTENNA__10876__A1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17815__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1143 _03417_ vssd1 vssd1 vccd1 vccd1 net2759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2770 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1165 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2781 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1176 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2792 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1187 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2803 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ net1088 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[4\] net907 vssd1
+ vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__and3_1
Xhold1198 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2814 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10628__A1 _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09494__A1 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08689_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[7\] net931 vssd1
+ vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10720_ _07058_ _07059_ net518 vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09121__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _06989_ _06990_ net537 vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10267__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15420__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10582_ net503 _06920_ vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__nand2_1
X_13370_ net1878 net826 _07650_ _03837_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12321_ net3252 net320 net434 vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__mux2_1
XANTENNA__12255__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10564__A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15040_ net1241 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__inv_2
XANTENNA__09549__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ net2814 net297 net442 vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__mux2_1
X_11203_ _06194_ _06218_ _07173_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__nand3_1
X_12183_ net3126 net299 net450 vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__mux2_1
XANTENNA__17345__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08969__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11134_ _07472_ _07473_ _07432_ vssd1 vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__a21o_1
X_18008__1508 vssd1 vssd1 vccd1 vccd1 _18008__1508/HI net1508 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_53_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16991_ clknet_leaf_7_wb_clk_i _02678_ _00974_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13502__B1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15942_ net1390 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__inv_2
X_11065_ _05454_ net374 _07371_ _07404_ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_120_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10016_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[1\] net738 _04687_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09721__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15873_ net1331 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14824_ net1289 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__inv_2
X_17612_ clknet_leaf_80_wb_clk_i _03297_ _01553_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17543_ clknet_leaf_124_wb_clk_i _03230_ _01526_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ net1350 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__inv_2
X_11967_ net3028 net275 net473 vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11334__S _07655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13706_ _04101_ _04123_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[3\]
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_47_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17474_ clknet_leaf_35_wb_clk_i _03161_ _01457_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10918_ _04738_ _06591_ _06917_ _05374_ _04736_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__a2111oi_1
X_17937__1437 vssd1 vssd1 vccd1 vccd1 _17937__1437/HI net1437 sky130_fd_sc_hd__conb_1
X_14686_ net1351 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11898_ net3127 net247 net480 vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16425_ clknet_leaf_104_wb_clk_i _02179_ _00408_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13637_ net200 net196 _07916_ net646 vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__o211a_1
X_10849_ _06469_ _06472_ _06568_ vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_15_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15330__A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16356_ clknet_leaf_78_wb_clk_i _02110_ _00339_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13568_ net197 net193 _07872_ net644 vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_97_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15307_ net1297 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12792__A1 _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12519_ net3087 net321 net410 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16287_ clknet_leaf_65_wb_clk_i net2613 _00270_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10474__A _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12165__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13499_ _03841_ _03951_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_93_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18026_ net1526 vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__buf_2
XFILLER_0_124_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15238_ net1292 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15169_ net1239 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__inv_2
Xfanout208 _07855_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16712__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09960__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout219 _07835_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__dlymetal6s2s_1
X_07991_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1 _04489_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_10_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09730_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[20\] net974
+ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_108_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_105_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10858__A1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09661_ _05999_ _06000_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__and2_1
XANTENNA__09206__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08612_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[11\] net652 net649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[11\]
+ _04951_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09592_ net512 vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09503__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08543_ net598 _04881_ _04882_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08474_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[23\] net907
+ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1070_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_A _07966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12783__A1 _07611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13980__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12075__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1335_A net1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09026_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[9\] net682 _05343_ _05349_
+ _05360_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_76_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout795_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold240 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold251 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[8\] vssd1 vssd1 vccd1 vccd1
+ net1878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 _01979_ vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold295 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[123\] vssd1 vssd1 vccd1 vccd1
+ net1911 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout962_A _04648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout720 net721 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_4
Xfanout731 net734 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_6
X_09928_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[4\] net819 net782 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__a22o_1
Xfanout742 _04685_ vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_8
Xfanout753 _04678_ vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__buf_6
XANTENNA__13496__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout764 net765 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_2
XANTENNA__08301__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout775 _04667_ vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__buf_6
Xfanout786 _04659_ vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__buf_6
Xfanout797 _04651_ vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__buf_4
X_09859_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[12\] _04634_ _04678_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[12\] vssd1 vssd1 vccd1 vccd1
+ _06199_ sky130_fd_sc_hd__a22o_1
XANTENNA__11510__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12870_ _04510_ _03575_ _03578_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_write_i
+ sky130_fd_sc_hd__nor3b_1
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11821_ net3169 net320 net494 vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14540_ net1392 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__inv_2
X_11752_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] _07938_ net615 vssd1
+ vssd1 vccd1 vccd1 _07939_ sky130_fd_sc_hd__mux2_4
XFILLER_0_16_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_132_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10703_ _07038_ _07042_ net528 vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14471_ net1333 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ net612 _07811_ _07883_ _07882_ vssd1 vssd1 vccd1 vccd1 _07884_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08690__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16210_ clknet_leaf_62_wb_clk_i net1752 _00198_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ _03861_ _03882_ _03860_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__a21oi_1
X_17190_ clknet_leaf_41_wb_clk_i _02877_ _01173_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12223__B1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10634_ _04707_ _05835_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_23_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12774__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16141_ clknet_leaf_95_wb_clk_i _01904_ _00129_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13353_ net566 _07678_ _03823_ _03825_ net586 vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__a32o_1
X_10565_ net531 net516 vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__nor2_2
XANTENNA__10785__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12304_ net1755 net239 net431 vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16072_ clknet_leaf_119_wb_clk_i _01865_ _00060_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_13284_ _04470_ _03752_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10496_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[31\] net942
+ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__and3_1
X_15023_ net1214 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12235_ net2703 net201 net439 vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__mux2_1
XANTENNA__12713__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10537__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12166_ net3136 net207 net447 vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11117_ _06921_ _07121_ vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__nor2_1
XANTENNA__12829__A2 _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ net3274 net247 net457 vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__mux2_1
X_16974_ clknet_leaf_6_wb_clk_i _02661_ _00957_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09155__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15925_ net1411 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__inv_2
X_11048_ _07386_ _07387_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__and2_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08363__D1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15325__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15856_ net1364 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16115__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08865__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14807_ net1195 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15787_ net1315 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12999_ net2327 net1805 net862 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14738_ net1318 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__inv_2
X_17526_ clknet_leaf_141_wb_clk_i _03213_ _01509_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08130__B2 _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11999__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17457_ clknet_leaf_15_wb_clk_i _03144_ _01440_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14669_ net1344 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__inv_2
XANTENNA__16265__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08881__B _05220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17510__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16408_ clknet_leaf_78_wb_clk_i _02162_ _00391_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08190_ net2351 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[83\] net1050 vssd1 vssd1
+ vccd1 vccd1 _03497_ sky130_fd_sc_hd__mux2_1
X_17388_ clknet_leaf_134_wb_clk_i _03075_ _01371_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12765__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16339_ clknet_leaf_86_wb_clk_i _02093_ _00322_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10240__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18009_ net1509 vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_hd__buf_2
XFILLER_0_23_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12623__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10528__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09933__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07974_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1 _04472_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09713_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[21\] net785 net753 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout376_A _05262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09644_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[23\] net821 net760 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09575_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[25\] net748 net741 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout543_A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1285_A net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08526_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[18\] net886 vssd1
+ vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_19_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11256__B2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08457_ net1084 net888 vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__and2_4
XANTENNA__17190__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18007__1507 vssd1 vssd1 vccd1 vccd1 _18007__1507/HI net1507 sky130_fd_sc_hd__conb_1
XANTENNA_fanout808_A net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16758__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08388_ net1156 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] _04624_ vssd1 vssd1
+ vccd1 vccd1 _04728_ sky130_fd_sc_hd__and3b_1
XFILLER_0_46_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12756__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10231__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[17\] net948
+ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12508__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[9\] net927 vssd1
+ vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10281_ _06608_ _06612_ _06616_ _06620_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__or4_1
XANTENNA__10519__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12533__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ net3202 net311 net468 vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11657__B net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__B _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17936__1436 vssd1 vssd1 vccd1 vccd1 _17936__1436/HI net1436 sky130_fd_sc_hd__conb_1
XFILLER_0_40_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16138__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout550 net552 vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__buf_2
XANTENNA__14130__B1 _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout561 _04749_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_4
Xfanout572 _04196_ vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__buf_1
X_13971_ _04218_ _04248_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__nor2_4
XFILLER_0_96_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout594 _04841_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_4
X_15710_ net1248 vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__inv_2
X_12922_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[16\] _03690_ net1032 vssd1
+ vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__mux2_1
X_16690_ clknet_leaf_129_wb_clk_i _02377_ _00673_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08685__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15641_ net1255 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__inv_2
X_12853_ net2509 net289 net381 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__mux2_1
XANTENNA__10289__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17533__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ net2530 net242 net491 vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__mux2_1
X_15572_ net1288 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08982__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12784_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] net1056 net365 _03617_
+ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17311_ clknet_leaf_24_wb_clk_i _02998_ _01294_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14523_ net1407 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11735_ _07922_ _07923_ _07925_ net613 vssd1 vssd1 vccd1 vccd1 _07926_ sky130_fd_sc_hd__a22o_4
XFILLER_0_132_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12708__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08663__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11612__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17242_ clknet_leaf_46_wb_clk_i _02929_ _01225_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14454_ net1369 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11666_ net2112 net241 net499 vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12747__A1 _07588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13405_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\]
+ net595 vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__and3_1
X_10617_ net541 _06953_ _06956_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17173_ clknet_leaf_123_wb_clk_i _02860_ _01156_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14385_ net1305 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__inv_2
Xwire940 _04756_ vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__clkbuf_2
X_11597_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _07813_ vssd1 vssd1
+ vccd1 vccd1 _07814_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16124_ clknet_leaf_109_wb_clk_i _01899_ _00112_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10222__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13336_ team_01_WB.instance_to_wrap.cpu.f0.i\[14\] _07681_ net564 vssd1 vssd1 vccd1
+ vccd1 _03812_ sky130_fd_sc_hd__o21ai_1
X_10548_ net508 _06098_ net543 vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16055_ clknet_leaf_92_wb_clk_i _01848_ _00043_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_126_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12443__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13267_ _03756_ _03758_ net2079 net829 vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__14224__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10479_ _06817_ _06818_ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15006_ net1274 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__inv_2
XANTENNA__09376__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ net3123 net311 net444 vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13198_ net10 net837 net630 net2080 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12149_ net1898 net279 net453 vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11286__C _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14121__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16957_ clknet_leaf_49_wb_clk_i _02644_ _00940_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11583__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15908_ net1398 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__inv_2
X_16888_ clknet_leaf_30_wb_clk_i _02575_ _00871_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09053__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15839_ net1372 vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11238__A1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09360_ _05687_ _05697_ _05698_ _05699_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__or4_1
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13632__C1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08311_ net989 net960 vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__and2_1
X_17509_ clknet_leaf_39_wb_clk_i _03196_ _01492_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16900__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09291_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[22\] net907 vssd1
+ vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__and3_1
XANTENNA__12618__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_126_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_13 _06589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08242_ net2837 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[31\] net1048 vssd1 vssd1
+ vccd1 vccd1 _03445_ sky130_fd_sc_hd__mux2_1
XANTENNA__10461__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_24 _07858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12738__A1 _07056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08173_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[108\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[100\]
+ net1039 vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__mux2_1
XANTENNA_68 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10213__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10764__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12353__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1033_A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_11_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09906__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XANTENNA__09228__A _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17406__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XANTENNA_fanout493_A _07944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput175 net175 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12910__A1 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1200_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14112__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07971__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16430__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17556__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08278__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09627_ _05965_ _05966_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout925_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09558_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] net626 _05897_ vssd1
+ vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__a21o_2
XFILLER_0_91_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08509_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[18\] net922
+ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10837__A net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[30\] net685 net655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__a22o_1
XANTENNA__12528__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11520_ team_01_WB.instance_to_wrap.cpu.DM0.enable net717 vssd1 vssd1 vccd1 vccd1
+ _07784_ sky130_fd_sc_hd__or2_2
XFILLER_0_68_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08307__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11451_ team_01_WB.instance_to_wrap.cpu.f0.i\[1\] _07671_ net327 vssd1 vssd1 vccd1
+ vccd1 _07750_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10275__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10402_ _06740_ _06741_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__nand2_1
X_14170_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\] _04189_ net1870 vssd1
+ vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11401__A1 _07696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13867__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11382_ _07710_ vssd1 vssd1 vccd1 vccd1 _07711_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09070__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13121_ net89 net845 net635 net2025 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a22o_1
XANTENNA__11668__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10333_ net559 _04883_ _05568_ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__or3_1
XANTENNA__12263__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09358__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ net2977 net2409 net859 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__mux2_1
XANTENNA_input54_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10264_ _06221_ _06603_ _06600_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__o21a_2
XFILLER_0_30_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12003_ net2305 net246 net467 vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__mux2_1
Xfanout1301 net1302 vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__clkbuf_4
X_10195_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[8\] net944 vssd1
+ vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1312 net1313 vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__buf_4
X_17860_ clknet_leaf_93_wb_clk_i _03535_ _01800_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.InstrRead
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1323 net1342 vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__clkbuf_8
Xfanout1334 net1335 vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08977__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14103__B1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1345 net1359 vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__clkbuf_2
X_16811_ clknet_leaf_5_wb_clk_i _02498_ _00794_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1356 net1358 vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__buf_4
X_17791_ clknet_leaf_62_wb_clk_i _03467_ _01731_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[61\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout1367 net1369 vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__buf_4
XFILLER_0_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout380 net382 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_6
Xfanout1378 net1379 vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__clkbuf_4
Xfanout1389 net1414 vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__buf_2
XANTENNA__11607__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout391 _03568_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_6
X_16742_ clknet_leaf_38_wb_clk_i _02429_ _00725_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13954_ _04217_ _04219_ _04222_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__and3_4
XANTENNA__08122__A2_N team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12905_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[21\] _03678_ net1031 vssd1
+ vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16673_ clknet_leaf_41_wb_clk_i _02360_ _00656_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13885_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[14\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[17\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_18_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13209__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15624_ net1277 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__inv_2
X_12836_ net2832 _07831_ net380 vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09601__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13090__A0 _03713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15555_ net1176 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10979__A0 _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[20\] _07171_ net1025 vssd1 vssd1
+ vccd1 vccd1 _03606_ sky130_fd_sc_hd__mux2_1
XANTENNA__12438__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14219__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14506_ net1387 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11718_ _07909_ _07911_ net612 vssd1 vssd1 vccd1 vccd1 _07912_ sky130_fd_sc_hd__mux2_8
X_15486_ net1248 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ net2998 net246 net383 vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__mux2_1
X_14437_ net1396 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__inv_2
X_17225_ clknet_leaf_9_wb_clk_i _02912_ _01208_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
X_11649_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] _07816_ vssd1 vssd1
+ vccd1 vccd1 _07857_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_1
XFILLER_0_109_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17156_ clknet_leaf_53_wb_clk_i _02843_ _01139_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput44 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16303__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14368_ net1343 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__inv_2
Xinput55 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput66 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
Xhold806 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[30\] vssd1 vssd1 vccd1 vccd1 net2422
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16107_ clknet_leaf_91_wb_clk_i _01882_ _00095_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold828 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ _07686_ _07706_ _03798_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] net586
+ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__o221a_1
XANTENNA__12173__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold839 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17087_ clknet_leaf_7_wb_clk_i _02774_ _01070_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14299_ net1352 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__inv_2
XANTENNA__09349__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09048__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16038_ clknet_leaf_103_wb_clk_i net1654 _00032_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08860_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[3\] net921 vssd1
+ vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18006__1506 vssd1 vssd1 vccd1 vccd1 _18006__1506/HI net1506 sky130_fd_sc_hd__conb_1
Xhold1506 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1517 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3133 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_106_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08791_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[0\] net896 vssd1
+ vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__and3_1
X_17989_ net1489 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
Xhold1528 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net3144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3155 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11517__S team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09521__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09412_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[27\] net679 net652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[27\]
+ _05741_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09343_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[25\] net899
+ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12348__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout241_A _07870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13620__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09230__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10434__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09274_ _05599_ _05602_ _05612_ _05613_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__or4_1
XFILLER_0_90_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08225_ net2717 net2691 net1049 vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1248_A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09588__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[125\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[117\]
+ net1040 vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10817__S0 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09884__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12083__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08087_ team_01_WB.instance_to_wrap.cpu.f0.i\[1\] _04524_ vssd1 vssd1 vccd1 vccd1
+ _04560_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout875_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16946__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[8\] net930 vssd1
+ vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09512__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ _06468_ _06471_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__nor2_1
XANTENNA__09124__C _04799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13670_ net1653 net567 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[31\] vssd1 vssd1
+ vccd1 vccd1 _01832_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10882_ _05566_ _06708_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12621_ _07791_ _07945_ net573 vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__and3_4
XFILLER_0_66_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08618__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15340_ net1206 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__inv_2
X_12552_ net2654 net319 net406 vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10425__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16326__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[11\] _07756_ vssd1 vssd1 vccd1
+ vccd1 _07779_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15271_ net1301 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__inv_2
X_12483_ net2362 net295 net414 vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17010_ clknet_leaf_130_wb_clk_i _02697_ _00993_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14222_ net1931 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09579__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13375__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11434_ _07676_ net610 _07737_ _04483_ _07699_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__a221oi_1
XANTENNA__10189__A1 _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14153_ _04416_ _04436_ net604 vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11365_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\] team_01_WB.instance_to_wrap.cpu.f0.i\[20\]
+ _07693_ vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13104_ net63 net62 _03726_ _03727_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__or4_1
X_10316_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[18\] net943
+ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__and3_1
X_14084_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[36\] _04221_ _04259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output160_A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11296_ net724 net644 vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13035_ net2368 net2091 net864 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__mux2_1
X_17912_ net1428 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
X_10247_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[9\] net784 net763 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[9\]
+ _06586_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__a221o_1
XANTENNA__14502__A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1120 net1121 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__clkbuf_2
Xfanout1131 net1132 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09751__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17843_ clknet_leaf_68_wb_clk_i net1681 _01783_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[113\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1142 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1 vccd1 vccd1
+ net1142 sky130_fd_sc_hd__buf_2
X_10178_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[10\] net740 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14088__C1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1153 net1154 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__clkbuf_2
Xfanout1164 net1167 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1175 net1177 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__buf_2
Xfanout1186 net1194 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__buf_4
X_17774_ clknet_leaf_56_wb_clk_i _03450_ _01714_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[44\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout1197 net1203 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__buf_4
X_14986_ net1272 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16725_ clknet_leaf_125_wb_clk_i _02412_ _00708_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13937_ _04227_ _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__nand2_4
XFILLER_0_92_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13868_ net1164 net1059 net1851 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[29\]
+ sky130_fd_sc_hd__and3b_1
X_16656_ clknet_leaf_126_wb_clk_i _02343_ _00639_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11580__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12819_ net1033 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[4\] vssd1 vssd1 vccd1
+ vccd1 _03642_ sky130_fd_sc_hd__or2_1
X_15607_ net1199 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12168__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13799_ _04170_ _04176_ _01838_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_100_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16587_ clknet_leaf_12_wb_clk_i _02274_ _00570_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_100_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13602__A2 _07553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15538_ net1233 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__inv_2
XANTENNA__17251__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15469_ net1208 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16819__CLK clknet_leaf_137_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08010_ team_01_WB.instance_to_wrap.a1.WRITE_I vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__inv_2
XANTENNA__11800__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17208_ clknet_leaf_27_wb_clk_i _02895_ _01191_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold603 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold614 _03432_ vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17139_ clknet_leaf_135_wb_clk_i _02826_ _01122_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold625 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold636 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 _02109_ vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09990__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09961_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[3\] net786 net745 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[3\]
+ _06292_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold669 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11129__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09209__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08912_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[2\] net684 _05232_ _05234_
+ _05238_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_102_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15508__A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09892_ net1134 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[5\] net968 vssd1
+ vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__and3_1
XANTENNA__12631__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08545__A1 net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ _05163_ _05164_ _05166_ _05168_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__or4_1
XFILLER_0_97_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09506__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1303 team_01_WB.instance_to_wrap.cpu.f0.num\[12\] vssd1 vssd1 vccd1 vccd1 net2919
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08410__A _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1314 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1325 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1336 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[14\] vssd1 vssd1 vccd1 vccd1
+ net2952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08774_ net599 _05110_ _05113_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__o21a_1
Xhold1347 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1358 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2974 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14094__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1369 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12867__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout456_A _07956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1198_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08783__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_74_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12078__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout623_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09326_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[24\] net698 net686 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09273__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09257_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[20\] net688 net668 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__a22o_1
XANTENNA__16499__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11080__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17744__CLK clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08208_ net2227 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[65\] net1050 vssd1 vssd1
+ vccd1 vccd1 _03479_ sky130_fd_sc_hd__mux2_1
XANTENNA__09025__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09188_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\] net703 _05510_ _05527_
+ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__o22a_4
XFILLER_0_62_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout992_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08139_ _04478_ team_01_WB.instance_to_wrap.cpu.f0.num\[16\] _04497_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\]
+ _04592_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a221o_1
XANTENNA__09981__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ _07476_ _07489_ vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__nor2_1
XANTENNA__09119__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10591__A1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ _06438_ _06440_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__and2_1
XANTENNA__12541__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ _07420_ _07353_ vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10032_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[0\] net941 vssd1
+ vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__and3_1
XANTENNA__09733__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14840_ net1179 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14085__A2 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ net1278 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__inv_2
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ net1818 net303 net472 vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__mux2_1
XANTENNA__13293__B1 _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08839__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16510_ clknet_leaf_112_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[8\]
+ _00493_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13722_ _04108_ _04130_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[12\]
+ sky130_fd_sc_hd__nor2_1
X_10934_ _05338_ net331 _07273_ net369 vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17490_ clknet_leaf_131_wb_clk_i _03177_ _01473_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17274__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16441_ clknet_leaf_39_wb_clk_i _02195_ _00424_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13653_ net188 _04085_ _04086_ net728 vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10865_ net339 _07201_ _07204_ net330 _07197_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12604_ net2712 net264 net395 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__mux2_1
XANTENNA__13596__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16372_ clknet_leaf_78_wb_clk_i _02126_ _00355_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13584_ _03900_ _03908_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__and2b_1
XANTENNA__08990__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09264__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10796_ _06036_ _07090_ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_45_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18111_ net636 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_45_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15323_ net1184 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__inv_2
X_18005__1505 vssd1 vssd1 vccd1 vccd1 _18005__1505/HI net1505 sky130_fd_sc_hd__conb_1
XFILLER_0_121_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12535_ net2099 net240 net403 vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12716__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18042_ net1542 vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15254_ net1201 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12466_ net3257 net201 net411 vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__mux2_1
X_14205_ net2775 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_1418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11417_ team_01_WB.instance_to_wrap.cpu.f0.i\[17\] _07690_ net325 vssd1 vssd1 vccd1
+ vccd1 _07732_ sky130_fd_sc_hd__o21ai_1
X_15185_ net1293 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__inv_2
X_12397_ net2740 net211 net420 vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08775__A1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14136_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[79\] _04235_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[119\]
+ _04420_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_91_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09972__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11348_ team_01_WB.instance_to_wrap.cpu.f0.i\[10\] team_01_WB.instance_to_wrap.cpu.f0.i\[9\]
+ net1064 vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__and3_2
XFILLER_0_39_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12451__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ net1169 _04329_ _04355_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10760__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14232__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ _07042_ _07099_ _07615_ _07618_ vssd1 vssd1 vccd1 vccd1 _07619_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13018_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[68\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[76\]
+ net856 vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__mux2_1
XANTENNA__11575__B _07784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10334__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11531__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17826_ clknet_leaf_75_wb_clk_i net1687 _01766_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14076__A2 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17757_ clknet_leaf_72_wb_clk_i net3051 _01697_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14969_ net1305 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11591__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10098__B1 _06436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16708_ clknet_leaf_50_wb_clk_i _02395_ _00691_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_08490_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[23\] net682 _04795_
+ _04807_ _04816_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10637__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17688_ clknet_leaf_94_wb_clk_i _03372_ _01629_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10919__B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15998__A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16639_ clknet_leaf_26_wb_clk_i _02326_ _00622_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09255__A2 _05591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09111_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[13\] net649 _05422_
+ _05430_ _05432_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_17_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12626__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wire960_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09042_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[12\] net917
+ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14000__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16791__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold400 _01966_ vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[12\] vssd1 vssd1 vccd1 vccd1 net2038
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A _07858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold433 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_121_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold444 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 net139 vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold466 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold477 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17147__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09944_ _06280_ _06283_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__and2_1
Xfanout902 net905 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__clkbuf_4
Xhold488 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 net916 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12361__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1113_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout924 _04767_ vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout935 net936 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13511__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08778__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout946 net947 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__buf_4
X_09875_ _06209_ _06213_ _06214_ net766 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__o32a_2
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout957 _04653_ vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__buf_4
Xhold1100 _02065_ vssd1 vssd1 vccd1 vccd1 net2716 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout968 _04640_ vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__clkbuf_8
Xhold1111 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[9\] vssd1 vssd1 vccd1 vccd1
+ net2727 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout979 _04629_ vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__buf_4
X_08826_ net1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[1\] net883 vssd1
+ vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_5_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1166 team_01_WB.instance_to_wrap.cpu.c0.count\[6\] vssd1 vssd1 vccd1 vccd1 net2782
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1177 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2793 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[4\] net892 vssd1
+ vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_87_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout740_A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1188 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1199 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[83\] vssd1 vssd1 vccd1 vccd1
+ net2815 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10089__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08688_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[7\] net888 vssd1
+ vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09494__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11006__A _05729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10650_ net512 _06811_ net548 vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__mux2_1
XANTENNA__09246__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09309_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[22\] net653 _05626_
+ _05640_ net706 vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_131_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10581_ _04710_ _06900_ vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__or2_4
XANTENNA__12536__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10845__A _06921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12320_ net2744 net306 net434 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08315__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10564__B _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ net2834 net299 net442 vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10013__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11202_ _07509_ _07520_ _07531_ _07541_ vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12182_ net2184 net282 net447 vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13367__S _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ _05189_ net331 _07433_ _06919_ net369 vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_129_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10580__A _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12271__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16990_ clknet_leaf_44_wb_clk_i _02677_ _00973_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_1450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13502__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16514__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08688__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15941_ net1411 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11064_ _05416_ net342 vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08914__D1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[1\] net804 net786 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__a22o_1
X_15872_ net1349 vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14058__A2 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08985__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17611_ clknet_leaf_80_wb_clk_i team_01_WB.instance_to_wrap.cpu.K0.next_keyvalid
+ _01552_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.keyvalid sky130_fd_sc_hd__dfrtp_4
X_14823_ net1299 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17542_ clknet_leaf_38_wb_clk_i _03229_ _01525_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11277__C1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14754_ net1315 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__inv_2
X_11966_ net2676 net211 net473 vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__mux2_1
XANTENNA__09485__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10917_ _05374_ _06591_ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__nand2_1
X_13705_ team_01_WB.instance_to_wrap.cpu.c0.count\[2\] team_01_WB.instance_to_wrap.cpu.c0.count\[1\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[0\] team_01_WB.instance_to_wrap.cpu.c0.count\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_47_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17473_ clknet_leaf_43_wb_clk_i _03160_ _01456_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14685_ net1344 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11897_ net3275 net213 net480 vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13569__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16424_ clknet_leaf_103_wb_clk_i _02178_ _00407_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13636_ _03862_ _03882_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__xnor2_1
X_10848_ net344 _07174_ _07175_ _07187_ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_89_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09237__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12938__A1_N _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12446__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16355_ clknet_leaf_86_wb_clk_i net2263 _00338_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_13567_ _03856_ _03920_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_97_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10779_ net530 _07118_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__nor2_1
XANTENNA__10755__A _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15306_ net1278 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12518_ net2224 net308 net410 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16286_ clknet_leaf_68_wb_clk_i _02040_ _00269_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13498_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] net981 _03957_ _03958_
+ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18025_ net1525 vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__buf_2
XANTENNA__16044__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12449_ net3223 net299 net417 vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__mux2_1
X_15237_ net1205 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__inv_2
X_15168_ net1242 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11752__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14119_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[6\] _04249_ _04262_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[54\]
+ _04398_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__a221o_1
XANTENNA__11586__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12181__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10490__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15099_ net1183 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__inv_2
X_07990_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1 _04488_
+ sky130_fd_sc_hd__inv_2
Xfanout209 net212 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_2
XANTENNA__16194__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09056__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09660_ net510 _05998_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10858__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14049__A2 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08611_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[11\] net902
+ net700 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[11\] vssd1 vssd1 vccd1
+ vccd1 _04951_ sky130_fd_sc_hd__a32o_1
X_17809_ clknet_leaf_77_wb_clk_i _03485_ _01749_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09591_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] net626 _05929_ _05930_
+ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__a22o_2
XFILLER_0_94_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08542_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] net619 net593 net600 vssd1
+ vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_82_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09476__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08473_ net1095 net906 vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_63_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout321_A _07937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10665__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12356__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout419_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09025_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[9\] net674 _05341_ _05352_
+ _05359_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_108_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1230_A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1328_A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09936__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07974__A team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold230 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[13\] vssd1 vssd1 vccd1 vccd1
+ net1846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold241 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[26\] vssd1 vssd1 vccd1 vccd1 net1857
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout690_A _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09892__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold252 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[23\] vssd1 vssd1 vccd1 vccd1
+ net1868 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[21\] vssd1 vssd1 vccd1 vccd1
+ net1890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold296 _02154_ vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout721 _04722_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_4
Xfanout732 net734 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09927_ _06257_ _06258_ _06259_ _06266_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_71_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_102_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout743 net745 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_6
Xfanout754 net755 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_8
Xfanout765 net767 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__buf_2
Xfanout776 _04667_ vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_6
Xfanout787 net788 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_8
X_09858_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[12\] net808 net787 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__a22o_1
X_18004__1504 vssd1 vssd1 vccd1 vccd1 _18004__1504/HI net1504 sky130_fd_sc_hd__conb_1
Xfanout798 net799 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__buf_6
XFILLER_0_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08809_ _05137_ _05140_ _05144_ _05148_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09789_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _06128_ net622 vssd1
+ vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__mux2_2
XFILLER_0_77_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11820_ net2094 net307 net494 vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11751_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[1\] _07476_ net718 vssd1 vssd1
+ vccd1 vccd1 _07938_ sky130_fd_sc_hd__mux2_1
XANTENNA__09132__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15431__A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10702_ _07039_ _07041_ net519 vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__mux2_1
XANTENNA__10278__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14470_ net1332 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _07809_ vssd1 vssd1
+ vccd1 vccd1 _07883_ sky130_fd_sc_hd__or2_1
XANTENNA__09219__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _03864_ _03881_ _03863_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10633_ net529 _06972_ _06966_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_23_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12266__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10234__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16140_ clknet_leaf_98_wb_clk_i _01903_ _00128_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12774__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13352_ _04486_ _07678_ _03824_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__o21a_1
XANTENNA__11431__C1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10564_ net558 _06902_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__or2_2
XANTENNA__10785__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ net3197 net271 net433 vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16071_ clknet_leaf_119_wb_clk_i _01864_ _00059_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_13283_ _04518_ _03747_ _03770_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__or3_1
XFILLER_0_126_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10495_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[31\] net811 vssd1 vssd1
+ vccd1 vccd1 _06835_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15022_ net1297 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__inv_2
X_12234_ net2304 net205 net439 vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17462__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12165_ net2137 net275 net448 vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ net525 _07200_ _07455_ vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_9_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12096_ net3264 net214 net457 vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__mux2_1
X_16973_ clknet_leaf_138_wb_clk_i _02660_ _00956_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09155__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11047_ net531 _06313_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__nand2_1
X_15924_ net1398 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12949__B net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09604__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15855_ net1364 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14806_ net1247 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15786_ net1315 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__inv_2
XANTENNA__09458__A2 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12998_ net2805 net2736 net860 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__mux2_1
XANTENNA__08666__A0 _04971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17525_ clknet_leaf_124_wb_clk_i _03212_ _01508_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09042__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14737_ net1320 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11949_ net2148 net302 net476 vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_116_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17456_ clknet_leaf_127_wb_clk_i _03143_ _01439_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14668_ net1355 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16407_ clknet_leaf_62_wb_clk_i _02161_ _00390_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12176__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13619_ _03888_ _04052_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17387_ clknet_leaf_5_wb_clk_i _03074_ _01370_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14599_ net1333 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16338_ clknet_leaf_61_wb_clk_i _02092_ _00321_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[61\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_27_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16269_ clknet_leaf_105_wb_clk_i net1743 _00257_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18008_ net1508 vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_hd__buf_2
XANTENNA__09918__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13190__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07973_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 _04471_
+ sky130_fd_sc_hd__inv_2
X_09712_ _06049_ _06050_ _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__or3_1
X_09643_ _05968_ _05981_ _05982_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__or3_1
XFILLER_0_39_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout369_A _06915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09574_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[25\] net947
+ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__and3_1
XANTENNA__09449__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08525_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[18\] net919 vssd1
+ vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__and3_1
XANTENNA__11256__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1180_A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1278_A net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08456_ net1112 net1114 net1107 net1110 vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__and4b_1
XANTENNA__07969__A team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_136_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09887__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08791__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12086__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08387_ _04626_ _04711_ net714 vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_46_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout703_A _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10767__A1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17485__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11003__B net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09008_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[9\] net911 vssd1
+ vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09909__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10280_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[19\] net731 _06617_ _06618_
+ _06619_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_44_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08312__B net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09127__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 _05189_ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__buf_2
Xfanout551 net552 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_4
Xfanout562 net563 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_4
X_13970_ _04218_ _04257_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__nor2_4
Xfanout573 _07961_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09688__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08966__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ _05528_ net577 net362 vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_57_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15640_ net1195 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__inv_2
X_12852_ net2622 net255 net379 vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ net3105 net273 net492 vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ net1281 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__inv_2
XANTENNA__11247__A2 _07524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12783_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[15\] _07611_ net1028 vssd1 vssd1
+ vccd1 vccd1 _03617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17310_ clknet_leaf_46_wb_clk_i _02997_ _01293_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10455__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14522_ net1394 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11734_ _07798_ _07924_ vssd1 vssd1 vccd1 vccd1 _07925_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09797__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09860__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16702__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17241_ clknet_leaf_55_wb_clk_i _02928_ _01224_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14453_ net1366 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__inv_2
X_11665_ _07867_ _07869_ net611 vssd1 vssd1 vccd1 vccd1 _07870_ sky130_fd_sc_hd__mux2_4
XANTENNA__10207__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10616_ net541 _06955_ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__nor2_1
X_13404_ _03863_ _03864_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__nand2b_1
X_14384_ net1305 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17172_ clknet_leaf_13_wb_clk_i _02859_ _01155_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11596_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\]
+ _07812_ vssd1 vssd1 vccd1 vccd1 _07813_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10758__A1 _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10758__B2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16123_ clknet_leaf_110_wb_clk_i _01898_ _00111_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13335_ _04480_ _07688_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__and2_1
X_10547_ _05837_ _06829_ _06885_ net344 vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__a31oi_1
XANTENNA__08820__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13266_ net825 _03757_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16054_ clknet_leaf_92_wb_clk_i _01847_ _00042_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_10478_ _06782_ _06814_ _06815_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11707__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13172__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12217_ net2241 net294 net446 vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__mux2_1
X_15005_ net1256 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__inv_2
X_13197_ net11 net837 net630 net2459 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12148_ net3276 net302 net453 vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09037__C _05374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10930__A1 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16956_ clknet_leaf_32_wb_clk_i _02643_ _00939_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08997__A2_N net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12079_ net3043 net228 net461 vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15907_ net1399 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__inv_2
XANTENNA__11583__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16887_ clknet_leaf_136_wb_clk_i _02574_ _00870_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16232__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08351__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17358__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15838_ net1358 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15769_ net1318 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11803__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08310_ net1147 net1149 net1152 net1154 vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__nor4b_2
X_17508_ clknet_leaf_55_wb_clk_i _03195_ _01491_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09290_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[22\] net889
+ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__and3_1
XANTENNA__16382__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10997__A1 _06915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10997__B2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08241_ net2560 net2456 net1046 vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_14 _06589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17439_ clknet_leaf_24_wb_clk_i _03126_ _01422_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09500__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 _07858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_36 _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_47 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[109\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[101\]
+ net1039 vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__mux2_1
XANTENNA_58 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_69 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18003__1503 vssd1 vssd1 vccd1 vccd1 _18003__1503/HI net1503 sky130_fd_sc_hd__conb_1
XANTENNA__08811__B1 _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12634__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_99_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09509__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08413__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
XANTENNA__09367__A1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13163__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_100_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XANTENNA__09228__B _05379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11174__A1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1026_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput176 net176 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08590__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08786__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout653_A _04819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1395_A net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09626_ _05963_ _05964_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09557_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\] net764 _05896_ net621
+ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout820_A _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08508_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[18\] net878
+ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09488_ _05820_ _05822_ _05827_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__or3_2
XANTENNA__09842__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08439_ net1114 net1112 net1109 net1106 vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__and4b_1
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11450_ _07673_ _07749_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ net372 _06739_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__or2_1
XANTENNA__12544__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ _04473_ _07709_ vssd1 vssd1 vccd1 vccd1 _07710_ sky130_fd_sc_hd__nor2_2
XFILLER_0_46_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ net90 net848 net631 net1825 vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10332_ _06671_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08323__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13051_ net2583 net2574 net864 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10263_ _06533_ _06594_ _06601_ _06602_ _06499_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__o32a_1
XFILLER_0_123_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10291__C net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ net2060 net201 net467 vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__mux2_1
Xfanout1302 net1303 vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__clkbuf_2
X_10194_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[8\] net802 net785 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input47_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10912__A1 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1313 net1314 vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__clkbuf_4
Xfanout1324 net1341 vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__buf_4
Xfanout1335 net1340 vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__buf_4
X_16810_ clknet_leaf_2_wb_clk_i _02497_ _00793_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1346 net1359 vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__buf_4
X_17790_ clknet_leaf_65_wb_clk_i _03466_ _01730_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[60\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__17500__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1357 net1358 vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__buf_4
Xfanout370 net371 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1368 net1369 vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__clkbuf_4
Xfanout381 net382 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_4
XANTENNA__09154__A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1379 net1380 vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__clkbuf_2
X_16741_ clknet_leaf_39_wb_clk_i _02428_ _00724_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout392 _03568_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_4
X_13953_ _04217_ _04220_ _04228_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__and3_4
XANTENNA__14995__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12904_ _05591_ net577 net361 vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_57_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16672_ clknet_leaf_29_wb_clk_i _02359_ _00655_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13884_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[11\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__or4bb_1
XANTENNA__08993__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10140__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15623_ net1301 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12417__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12835_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[30\] net223 net379 vssd1
+ vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12719__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10428__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11623__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15554_ net1266 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12766_ net1848 net639 net609 _03605_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10979__A1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09833__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14505_ net1398 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__inv_2
X_11717_ _07801_ _07910_ vssd1 vssd1 vccd1 vccd1 _07911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12697_ net2847 net203 net383 vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__mux2_1
X_15485_ net1263 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17224_ clknet_leaf_23_wb_clk_i _02911_ _01207_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14436_ net1400 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__inv_2
X_11648_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[22\] _07154_ net715 vssd1 vssd1
+ vccd1 vccd1 _07856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 gpio_in[16] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_1
XFILLER_0_29_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17155_ clknet_leaf_19_wb_clk_i _02842_ _01138_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput45 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12454__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14367_ net1343 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__inv_2
X_11579_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[31\] _06961_ net715 vssd1 vssd1
+ vccd1 vccd1 _07796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput56 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_1
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold807 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[97\] vssd1 vssd1 vccd1 vccd1
+ net2423 sky130_fd_sc_hd__dlygate4sd3_1
Xinput67 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dlymetal6s2s_1
X_16106_ clknet_leaf_91_wb_clk_i _01881_ _00094_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13318_ team_01_WB.instance_to_wrap.cpu.f0.i\[17\] net610 _07703_ vssd1 vssd1 vccd1
+ vccd1 _03798_ sky130_fd_sc_hd__and3_1
Xhold818 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
X_17086_ clknet_leaf_45_wb_clk_i _02773_ _01069_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold829 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[78\] vssd1 vssd1 vccd1 vccd1
+ net2445 sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ net1352 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__inv_2
XANTENNA__13145__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16037_ clknet_leaf_103_wb_clk_i _01831_ _00031_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13249_ net2312 net356 net352 team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1
+ vccd1 vccd1 _01901_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11594__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17180__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1507 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3123 sky130_fd_sc_hd__dlygate4sd3_1
X_08790_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[0\] net925 vssd1
+ vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17988_ net1488 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
Xhold1518 team_01_WB.instance_to_wrap.cpu.f0.num\[28\] vssd1 vssd1 vccd1 vccd1 net3134
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3145 sky130_fd_sc_hd__dlygate4sd3_1
X_16939_ clknet_leaf_4_wb_clk_i _02626_ _00922_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09411_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[27\] net683 _05750_
+ net707 vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__a211o_1
XANTENNA__12629__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16898__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ _05681_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__inv_2
XANTENNA__12959__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08088__B2 team_01_WB.instance_to_wrap.cpu.f0.write_data\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08408__A _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09273_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[20\] net651 net649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[20\]
+ _05598_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout234_A _07884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08224_ net2068 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[49\] net1050 vssd1 vssd1
+ vccd1 vccd1 _03463_ sky130_fd_sc_hd__mux2_1
XANTENNA__10376__C net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14030__B1 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08155_ net1786 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[118\] net1042 vssd1 vssd1
+ vccd1 vccd1 _03532_ sky130_fd_sc_hd__mux2_1
XANTENNA__12364__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout401_A _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10817__S1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1143_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08086_ _04529_ _04539_ _04558_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_3_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1408_A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13541__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout770_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout868_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14097__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[8\] net935 vssd1
+ vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10658__A0 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__A _05707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ net563 _07189_ _07270_ _07289_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__a31o_2
XANTENNA__10122__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09609_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[24\] net783 net773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__a22o_1
X_10881_ _05566_ net331 _07220_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12539__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12620_ net2151 net291 net396 vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09276__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09815__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12551_ net2122 net307 net405 vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__mux2_1
XANTENNA__11083__B1 _05707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ net1657 net876 _07758_ _07778_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__o22a_1
X_12482_ net2389 net299 net414 vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17053__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15270_ net1290 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14021__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14221_ net2082 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13375__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11433_ _07678_ _07701_ _07741_ net326 vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__o211a_1
XANTENNA__12274__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14055__A _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14152_ _04222_ _04228_ _04237_ _04289_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__a31o_1
X_11364_ team_01_WB.instance_to_wrap.cpu.f0.i\[19\] _07692_ vssd1 vssd1 vccd1 vccd1
+ _07693_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10315_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[18\] net969 vssd1
+ vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__and3_1
X_13103_ net59 net60 vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14083_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[60\] _04260_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[116\]
+ _04370_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11295_ net726 _04838_ vssd1 vssd1 vccd1 vccd1 _07635_ sky130_fd_sc_hd__nor2_1
XANTENNA__08988__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13034_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[52\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[60\]
+ net856 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__mux2_1
X_17911_ net1427 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
X_10246_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[9\] _04654_ _06584_
+ _06585_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12886__A1 _05726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1110 net1111 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11618__S net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1121 net1127 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__buf_2
X_17842_ clknet_leaf_75_wb_clk_i net2532 _01782_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[112\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1132 net1135 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__buf_2
X_10177_ _06505_ _06508_ _06513_ _06516_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__nor4_1
Xfanout1143 net1145 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__buf_2
Xfanout1154 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] vssd1 vssd1 vccd1 vccd1
+ net1154 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1165 net1166 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__clkbuf_2
Xfanout1176 net1177 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__buf_4
X_17773_ clknet_leaf_72_wb_clk_i net3242 _01713_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_18079__1579 vssd1 vssd1 vccd1 vccd1 _18079__1579/HI net1579 sky130_fd_sc_hd__conb_1
X_14985_ net1229 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__inv_2
Xfanout1187 net1194 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__clkbuf_4
Xfanout1198 net1203 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__clkbuf_4
X_18002__1502 vssd1 vssd1 vccd1 vccd1 _18002__1502/HI net1502 sky130_fd_sc_hd__conb_1
XFILLER_0_135_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10649__A0 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16724_ clknet_leaf_12_wb_clk_i _02411_ _00707_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13936_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__nor2_4
XFILLER_0_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11310__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16655_ clknet_leaf_144_wb_clk_i _02342_ _00638_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12449__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13867_ net1164 net1059 net1697 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[28\]
+ sky130_fd_sc_hd__and3b_1
X_15606_ net1247 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__inv_2
X_12818_ net1034 _07449_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__nand2_1
XANTENNA__11580__C team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09267__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16586_ clknet_leaf_11_wb_clk_i _02273_ _00569_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_13798_ _04159_ _04174_ _04179_ _04154_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09806__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15537_ net1341 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__inv_2
XANTENNA__09050__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12749_ net1919 net639 net606 _03593_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a22o_1
XANTENNA__11613__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12810__B2 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10196__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14012__B1 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15468_ net1205 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17207_ clknet_leaf_140_wb_clk_i _02894_ _01190_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14419_ net1366 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12184__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16420__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15399_ net1328 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13771__C1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09059__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17138_ clknet_leaf_129_wb_clk_i _02825_ _01121_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold604 team_01_WB.instance_to_wrap.cpu.f0.state\[7\] vssd1 vssd1 vccd1 vccd1 net2220
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold615 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold626 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold637 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09960_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[3\] net748 net737 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__a22o_1
X_17069_ clknet_leaf_140_wb_clk_i _02756_ _01052_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08898__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13523__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08911_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[2\] net681 _05230_ _05236_
+ _05240_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17696__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09891_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[5\] _04665_
+ vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12877__A1 _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08545__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08842_ _05179_ _05180_ _05181_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__or3_1
XANTENNA__14079__B1 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1304 _01912_ vssd1 vssd1 vccd1 vccd1 net2920 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08410__B net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10352__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1315 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1326 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[119\] vssd1 vssd1 vccd1 vccd1
+ net2942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08773_ net602 _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__or2_1
Xhold1337 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1348 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1359 team_01_WB.instance_to_wrap.cpu.c0.count\[4\] vssd1 vssd1 vccd1 vccd1 net2975
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12359__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1093_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_A _07958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_942 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09258__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17076__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09325_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[24\] net679 net672 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[24\]
+ _05663_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12801__A1 _07269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1260_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1358_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[20\] net933
+ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14003__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08207_ net2624 net2437 net1043 vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_43_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09187_ _05514_ _05518_ _05522_ _05526_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12094__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08138_ _04478_ team_01_WB.instance_to_wrap.cpu.f0.num\[16\] team_01_WB.instance_to_wrap.cpu.f0.num\[10\]
+ _04483_ _04591_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_47_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09430__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout985_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16913__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08784__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08304__C net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__B net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08069_ _04542_ _04543_ _04544_ _04545_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10100_ _05043_ _06439_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11080_ _05618_ net507 _07355_ net508 _05594_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__o32a_1
XFILLER_0_80_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10031_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[0\] net947 vssd1
+ vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__and3_1
XANTENNA__08536__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11540__B2 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09135__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14770_ net1326 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ net2250 net284 net473 vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__mux2_1
XANTENNA__08974__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17419__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13721_ net2267 _04107_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__nor2_1
X_10933_ _06919_ net336 _07272_ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12269__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16440_ clknet_leaf_20_wb_clk_i _02194_ _00423_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10864_ _07118_ _07200_ net525 vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__mux2_1
X_13652_ net200 net196 _07930_ net646 vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__o211a_1
XANTENNA__09249__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13889__A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12603_ net2393 net270 net395 vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16371_ clknet_leaf_85_wb_clk_i _02125_ _00354_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13596__A2 _07188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16443__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10795_ net562 _07115_ _07116_ _07134_ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__a31o_2
X_13583_ net984 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] _04027_ _04028_
+ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a22o_1
XANTENNA__17569__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18110_ net636 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11901__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15322_ net1189 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__inv_2
X_12534_ net3142 net273 net405 vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18041_ net1541 vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__buf_2
X_15253_ net1222 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12465_ net3239 net205 net411 vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14204_ net3019 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_1532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11416_ _07692_ net325 _07730_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__and3b_1
XFILLER_0_105_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15184_ net1270 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__inv_2
X_12396_ net1950 net248 net422 vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09421__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14135_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[87\] _04251_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[79\]
+ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__a22o_1
XANTENNA__08775__A2 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11347_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\] _07675_ vssd1 vssd1 vccd1 vccd1
+ _07676_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_91_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09607__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12859__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14066_ _04332_ _04341_ _04348_ _04354_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__or4_1
X_11278_ _05595_ net508 _07616_ _07617_ vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__o22a_1
XANTENNA__08511__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09724__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13017_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[69\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[77\]
+ net855 vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__mux2_1
X_10229_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[9\] net776 _04678_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__a22o_1
XANTENNA__11575__C _07789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11531__B2 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17825_ clknet_leaf_77_wb_clk_i net3187 _01765_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1 team_01_WB.instance_to_wrap.cpu.K0.state vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09045__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17756_ clknet_leaf_66_wb_clk_i net2230 _01696_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_76_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14968_ net1178 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10098__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16707_ clknet_leaf_23_wb_clk_i _02394_ _00690_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11591__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13919_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\] _04212_ _04213_ vssd1
+ vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__o21a_1
XANTENNA__12179__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17687_ clknet_leaf_96_wb_clk_i _03371_ _01628_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14899_ net1234 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16638_ clknet_leaf_44_wb_clk_i _02325_ _00621_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16569_ clknet_leaf_58_wb_clk_i _02256_ _00552_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09110_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[13\] net684 _05421_
+ _05442_ net709 vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11811__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16936__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09041_ net1155 net619 net593 vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold401 net91 vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09412__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold412 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold434 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12642__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold445 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold456 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[6\] vssd1 vssd1 vccd1 vccd1
+ net2072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11770__A1 _07866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold478 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09943_ _05115_ _06282_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__xnor2_1
Xhold489 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[31\] vssd1 vssd1 vccd1 vccd1
+ net2105 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout903 net904 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__buf_4
XANTENNA__10670__B _06398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout914 net916 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout925 net926 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__buf_4
XANTENNA__10493__A_N net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout936 _04759_ vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout399_A _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13511__A2 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[12\] net751 net749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[12\]
+ _06197_ vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__a221o_1
Xfanout947 _04662_ vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_8
Xfanout958 _04653_ vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_4
Xhold1101 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[56\] vssd1 vssd1 vccd1 vccd1
+ net2717 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16316__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11522__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout969 _04638_ vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__clkbuf_8
Xhold1112 _02048_ vssd1 vssd1 vccd1 vccd1 net2728 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[1\] net908 vssd1
+ vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__and3_1
Xhold1123 team_01_WB.instance_to_wrap.cpu.f0.num\[8\] vssd1 vssd1 vccd1 vccd1 net2739
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1134 team_01_WB.instance_to_wrap.cpu.f0.num\[5\] vssd1 vssd1 vccd1 vccd1 net2750
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2772 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1167 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08756_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[4\] net923 vssd1
+ vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_87_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1178 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2794 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13275__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[88\] vssd1 vssd1 vccd1 vccd1
+ net2805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12089__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout733_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08687_ net1073 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[7\] net938 vssd1
+ vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout900_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09308_ _05644_ _05645_ _05646_ _05647_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__or4_1
X_10580_ _04710_ _06900_ vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_131_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09651__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09239_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[21\] net688 net666 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_40_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18078__1578 vssd1 vssd1 vccd1 vccd1 _18078__1578/HI net1578 sky130_fd_sc_hd__conb_1
XFILLER_0_44_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12250_ net3073 net279 net439 vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__mux2_1
X_18001__1501 vssd1 vssd1 vccd1 vccd1 _18001__1501/HI net1501 sky130_fd_sc_hd__conb_1
XANTENNA__09403__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11201_ _07533_ _07539_ _07540_ vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__or3_4
X_12181_ net2020 net304 net449 vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__mux2_1
XANTENNA__12552__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ net338 _07433_ vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_129_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08969__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11063_ _07379_ _07402_ vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__nand2_1
X_15940_ net1388 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__inv_2
XANTENNA__13502__A2 _07019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10014_ _06350_ _06351_ _06352_ _06353_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_34_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09182__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15871_ net1347 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__inv_2
X_17610_ clknet_leaf_80_wb_clk_i team_01_WB.instance_to_wrap.cpu.K0.next_state _01551_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.state sky130_fd_sc_hd__dfrtp_1
X_14822_ net1299 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__inv_2
XANTENNA__09162__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17541_ clknet_leaf_38_wb_clk_i _03228_ _01524_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14753_ net1316 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11965_ net2289 net249 net473 vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13704_ net2975 _04101_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[4\]
+ sky130_fd_sc_hd__xor2_1
X_17472_ clknet_leaf_30_wb_clk_i _03159_ _01455_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10916_ _07254_ _07255_ net519 vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10101__A _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_106_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14684_ net1348 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__inv_2
X_11896_ net2930 net219 net479 vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16959__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16423_ clknet_leaf_104_wb_clk_i _02177_ _00406_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ net982 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] _04071_ _04072_
+ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ net554 _07186_ _07184_ vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_32_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11631__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16354_ clknet_leaf_61_wb_clk_i _02108_ _00337_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[77\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_15_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13566_ net980 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] _04013_ _04014_
+ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10778_ _07104_ _07117_ net514 vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10755__B net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15305_ net1230 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__inv_2
XANTENNA__10252__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12517_ net2853 net310 net408 vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16285_ clknet_leaf_84_wb_clk_i net2411 _00268_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13497_ net724 _06961_ net1067 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_93_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18024_ net1524 vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__buf_2
X_15236_ net1191 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12448_ net2341 net281 net415 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12462__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15167_ net1255 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__inv_2
X_12379_ net2203 net253 net425 vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__mux2_1
XANTENNA__14243__A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14118_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[46\] _04246_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[126\]
+ _04403_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11586__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15098_ net1190 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14151__C1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14049_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[91\] _04241_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[59\]
+ _04337_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10858__A3 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_4__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11806__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08920__A2 _05258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[11\] net688 net653 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__a22o_1
XANTENNA__15074__A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17808_ clknet_leaf_65_wb_clk_i net2910 _01748_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_09590_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\] net765 net622 vssd1
+ vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__o21a_1
XANTENNA__17734__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17739_ clknet_leaf_71_wb_clk_i _03415_ _01679_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_08541_ net592 net591 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] net702
+ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__o2bb2a_4
XTAP_TAPCELL_ROW_82_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09503__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08472_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[23\] net878
+ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__and3_1
XANTENNA__15802__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12733__B1_N net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17884__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12637__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13322__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08987__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13980__A2 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17114__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout314_A _07939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[9\] net671 _05345_ _05351_
+ _05354_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1056_A team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13193__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 _01983_ vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12372__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold231 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[24\] vssd1 vssd1 vccd1 vccd1
+ net1847 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1223_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold242 _01992_ vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12940__B1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08789__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold264 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 _04760_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__buf_6
Xhold286 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout683_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold297 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[121\] vssd1 vssd1 vccd1 vccd1
+ net1913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09926_ _06260_ _06261_ _06265_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__or3_1
Xfanout722 net724 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__clkbuf_4
Xfanout733 net734 vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_6
XANTENNA__13496__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout744 net745 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_4
Xfanout755 _04676_ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__buf_6
XANTENNA__07990__A team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout766 net767 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout777 net778 vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_8
X_09857_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[12\] net965
+ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout850_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout788 _04657_ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout799 _04649_ vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout948_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08911__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08808_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[0\] net685 _05145_ _05146_
+ _05147_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13248__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09788_ _06111_ _06118_ _06126_ _06127_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__o31a_1
X_08739_ net1008 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[4\] net930 vssd1
+ vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ net3269 net320 net502 vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09872__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10701_ _07040_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11681_ net720 _07611_ net615 _07881_ vssd1 vssd1 vccd1 vccd1 _07882_ sky130_fd_sc_hd__o211a_1
XANTENNA__12547__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _03867_ _03880_ _03866_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ net515 _06969_ _06970_ _06971_ vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_23_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10563_ net558 _06902_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13351_ team_01_WB.instance_to_wrap.cpu.f0.i\[11\] _07685_ vssd1 vssd1 vccd1 vccd1
+ _03824_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10785__A2 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12302_ net3236 net243 net431 vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16070_ clknet_leaf_120_wb_clk_i _01863_ _00058_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\]
+ sky130_fd_sc_hd__dfstp_4
X_10494_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[31\] net978
+ vssd1 vssd1 vccd1 vccd1 _06834_ sky130_fd_sc_hd__and3_1
X_13282_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] _03746_ team_01_WB.instance_to_wrap.cpu.f0.i\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15021_ net1207 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__inv_2
XANTENNA__13184__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11687__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12282__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12233_ net3056 net276 net441 vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10537__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12931__B1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09157__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12164_ net2287 net211 net448 vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11115_ _06905_ _07303_ _07454_ _05263_ vssd1 vssd1 vccd1 vccd1 _07455_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_124_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16972_ clknet_leaf_133_wb_clk_i _02659_ _00955_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16631__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12095_ net2981 net219 net457 vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_55_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11046_ net531 _06313_ vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__or2_1
X_15923_ net1402 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__inv_2
XANTENNA__09155__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11626__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15854_ net1364 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__inv_2
XANTENNA__10170__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13239__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_95_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16781__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14805_ net1220 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__inv_2
X_15785_ net1309 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__inv_2
X_12997_ net2856 net2830 net867 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17524_ clknet_leaf_12_wb_clk_i _03211_ _01507_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14736_ net1320 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__inv_2
X_11948_ net2191 net283 net477 vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__mux2_1
XANTENNA__08666__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ clknet_leaf_143_wb_clk_i _03142_ _01438_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12457__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14667_ net1376 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__inv_2
X_11879_ net2479 net289 net486 vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16406_ clknet_leaf_62_wb_clk_i _02160_ _00389_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13618_ net982 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] _04057_ _04058_
+ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17386_ clknet_leaf_10_wb_clk_i _03073_ _01369_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14598_ net1334 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16337_ clknet_leaf_64_wb_clk_i _02091_ _00320_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[60\]
+ sky130_fd_sc_hd__dfstp_1
X_13549_ net980 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] _03999_ _04000_
+ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16268_ clknet_leaf_105_wb_clk_i net1733 _00256_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
XANTENNA__17287__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18007_ net1507 vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_hd__buf_2
XANTENNA__13175__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15219_ net1280 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11597__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12192__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16199_ clknet_leaf_114_wb_clk_i _01959_ _00187_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10528__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07972_ team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 _04470_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09711_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[21\] net760 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08354__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09642_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[23\] net807 _05972_
+ _05974_ _05980_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_39_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18077__1577 vssd1 vssd1 vccd1 vccd1 _18077__1577/HI net1577 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_65_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09573_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[25\] net942
+ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__and3_1
X_18000__1500 vssd1 vssd1 vccd1 vccd1 _18000__1500/HI net1500 sky130_fd_sc_hd__conb_1
XANTENNA__08106__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08524_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[18\] net897 vssd1
+ vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09530__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08455_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[23\] net893 vssd1
+ vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__and3_1
XANTENNA__12367__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1173_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08386_ net1156 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\] _04623_ _04725_ vssd1
+ vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_78_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1340_A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13166__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout898_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09007_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[9\] net884 vssd1
+ vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__and3_1
XANTENNA__09909__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16654__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10519__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09385__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout530 net532 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_2
Xfanout541 net542 vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_4
X_09909_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\] net766 net623 vssd1
+ vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__o21a_1
XANTENNA__14130__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout552 _05151_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_2
XANTENNA__09705__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout563 _04747_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_4
Xfanout574 _07961_ vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_1
Xfanout585 net586 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__buf_2
XFILLER_0_77_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12920_ net358 _03688_ _03689_ net871 net2212 vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a32o_1
Xfanout596 net597 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10152__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12851_ net3013 net260 net382 vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_9__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_48_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13626__D1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10289__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15442__A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[21\] net243 net491 vssd1
+ vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ net1234 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12782_ net1712 net641 net608 _03616_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08982__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14521_ net1398 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11733_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] _07797_ vssd1 vssd1 vccd1
+ vccd1 _07924_ sky130_fd_sc_hd__nor2_1
XANTENNA__12277__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17240_ clknet_leaf_25_wb_clk_i _02927_ _01223_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14452_ net1368 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__inv_2
XANTENNA__16184__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11664_ _07813_ _07868_ vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] net596 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__a21o_1
X_10615_ net547 _06366_ _06399_ vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17171_ clknet_leaf_128_wb_clk_i _02858_ _01154_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14383_ net1308 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__inv_2
X_11595_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\]
+ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _07809_ vssd1 vssd1 vccd1 vccd1
+ _07812_ sky130_fd_sc_hd__and4_1
XFILLER_0_51_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10758__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16122_ clknet_leaf_100_wb_clk_i _01897_ _00110_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13334_ net2469 net829 _03809_ _03810_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__a22o_1
X_10546_ _05837_ _06829_ _06885_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13157__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16053_ clknet_leaf_92_wb_clk_i _01846_ _00041_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_13265_ _04518_ _03750_ _03755_ _04621_ _04466_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__o221ai_1
X_10477_ net512 _05933_ _06816_ vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__o21ai_2
XANTENNA__11707__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15004_ net1172 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__inv_2
X_12216_ net2605 net300 net446 vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09376__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13196_ net12 net837 net630 net2551 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_63_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12147_ net2120 net283 net452 vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10391__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10930__A2 _06472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14121__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16955_ clknet_leaf_20_wb_clk_i _02642_ _00938_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12078_ net2032 net287 net461 vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__mux2_1
X_15906_ net1383 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__inv_2
X_11029_ _05455_ net374 vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__nor2_1
XANTENNA__10143__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16886_ clknet_leaf_141_wb_clk_i _02573_ _00869_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15837_ net1372 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__inv_2
XANTENNA__09053__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10199__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15768_ net1321 vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09836__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13632__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16527__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08892__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17507_ clknet_leaf_23_wb_clk_i _03194_ _01490_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14719_ net1315 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12187__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15699_ net1280 vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__inv_2
XANTENNA__10496__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08240_ net2023 net2587 net1050 vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__mux2_1
X_17438_ clknet_leaf_44_wb_clk_i _03125_ _01421_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_15 _06737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_26 _07858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08171_ net2821 net2592 net1044 vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__mux2_1
XANTENNA_48 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17369_ clknet_leaf_51_wb_clk_i _03056_ _01352_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16677__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_59 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08811__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13148__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_113_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_105_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_81_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XFILLER_0_100_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_0_10_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput177 net177 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XANTENNA__12650__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10382__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14112__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout381_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12123__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13850__A_N net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13320__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A _07949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17302__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09625_ _05963_ _05964_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1290_A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1388_A net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09556_ _05888_ _05889_ _05893_ _05895_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__or4_2
XANTENNA__09827__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13623__A1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17452__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08507_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] net619 net593 vssd1 vssd1
+ vccd1 vccd1 _04847_ sky130_fd_sc_hd__a21o_1
XANTENNA__12097__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11634__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ _05823_ _05824_ _05825_ _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout813_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08438_ net1010 net930 vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__and2_4
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08307__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11014__B net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08369_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] net1155 vssd1 vssd1 vccd1
+ vccd1 _04709_ sky130_fd_sc_hd__and2b_1
XFILLER_0_92_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11937__A1 _07866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10400_ net372 _06739_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__nand2_2
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11380_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] _07707_ vssd1 vssd1 vccd1 vccd1
+ _07709_ sky130_fd_sc_hd__nand2_2
XANTENNA__13139__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10331_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] net625 _06669_ _06670_
+ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__a22o_4
XFILLER_0_132_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08323__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13050_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[36\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[44\]
+ net855 vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__mux2_1
X_10262_ _06500_ _06530_ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__nor2_1
XANTENNA__09358__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09138__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ net2406 net205 net467 vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__mux2_1
X_10193_ _06499_ _06500_ _06532_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__or3_1
XANTENNA__12560__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1303 net1415 vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__buf_2
Xfanout1314 net1342 vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__buf_2
Xfanout1325 net1329 vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__buf_4
XANTENNA__10912__A2 _06472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14103__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08977__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1336 net1340 vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__buf_4
Xfanout1347 net1359 vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__buf_2
Xfanout360 _03655_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1358 net1359 vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout371 _06914_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13311__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1369 net1380 vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__buf_2
X_16740_ clknet_leaf_50_wb_clk_i _02427_ _00723_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout382 _03651_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_8
X_13952_ _04220_ _04237_ _04239_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__and3_4
Xfanout393 _03568_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_8
XANTENNA__10125__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10676__A1 _07015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12903_ net358 _03676_ _03677_ net871 net2548 vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__a32o_1
X_16671_ clknet_leaf_26_wb_clk_i _02358_ _00654_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13883_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[7\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__or4b_1
XFILLER_0_92_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11904__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15622_ net1296 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__inv_2
XANTENNA__09818__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12834_ net2620 net190 net380 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15553_ net1250 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__inv_2
X_12765_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] net1054 net364 _03604_
+ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__a22o_1
XANTENNA__09601__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10979__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14504_ net1384 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11716_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] _07800_ vssd1 vssd1 vccd1
+ vccd1 _07910_ sky130_fd_sc_hd__nor2_1
X_15484_ net1171 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12696_ net2894 net205 net383 vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17223_ clknet_leaf_16_wb_clk_i _02910_ _01206_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14435_ net1396 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__inv_2
X_11647_ net3040 net207 net499 vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_1
XFILLER_0_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17154_ clknet_leaf_36_wb_clk_i _02841_ _01137_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput35 gpio_in[17] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
XFILLER_0_13_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14366_ net1349 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11578_ net576 _07793_ _07794_ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__and3_4
XANTENNA__08514__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput46 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
Xinput57 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput68 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
X_16105_ clknet_leaf_91_wb_clk_i _01880_ _00093_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18076__1576 vssd1 vssd1 vccd1 vccd1 _18076__1576/HI net1576 sky130_fd_sc_hd__conb_1
Xhold808 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 net2424
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13317_ net1975 net825 _03795_ _03797_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__o22a_1
XFILLER_0_40_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17085_ clknet_leaf_21_wb_clk_i _02772_ _01068_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold819 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[79\] vssd1 vssd1 vccd1 vccd1
+ net2435 sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[31\] net676 net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[31\]
+ _06868_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__a221o_1
X_14297_ net1355 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16036_ clknet_leaf_102_wb_clk_i _01830_ _00030_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09349__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13248_ net2734 net355 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1
+ vccd1 vccd1 _01902_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09048__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15347__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17325__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12470__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ net1671 net851 net841 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_1203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08887__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09345__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11594__B _07809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1508 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3124 sky130_fd_sc_hd__dlygate4sd3_1
X_17987_ net1487 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
Xhold1519 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16938_ clknet_leaf_3_wb_clk_i _02625_ _00921_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09521__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16869_ clknet_leaf_38_wb_clk_i _02556_ _00852_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11814__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[27\] net695 _04808_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[27\] vssd1 vssd1 vccd1 vccd1
+ _05750_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09341_ net599 _05678_ _05680_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09272_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[20\] net683 _05611_
+ net707 vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_115_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13369__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08223_ net2616 net2481 net1043 vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12645__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout227_A _07900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08154_ net1709 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[119\] net1046 vssd1 vssd1
+ vccd1 vccd1 _03533_ sky130_fd_sc_hd__mux2_1
XANTENNA__09588__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08085_ _04515_ _04523_ _04537_ _04557_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout1136_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout596_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1303_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12895__A2 _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[8\] net662 _05325_ _05326_
+ net709 vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__17818__CLK clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout763_A _04674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10107__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10658__A1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11009__B net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout930_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08720__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09608_ net992 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[24\] net976 vssd1
+ vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16842__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10880_ _05566_ _06708_ net369 vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[28\] net962
+ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__and3_1
XANTENNA__09276__A1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15720__A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12550_ net2958 net313 net404 vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__mux2_1
XANTENNA__11083__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16992__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11501_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[12\] _07756_ vssd1 vssd1 vccd1
+ vccd1 _07778_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ net2408 net279 net411 vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14220_ net2188 vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__clkbuf_1
X_11432_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\] _07675_ net610 team_01_WB.instance_to_wrap.cpu.f0.i\[11\]
+ vssd1 vssd1 vccd1 vccd1 _07741_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09579__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08334__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14055__B _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12583__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14151_ net1761 net604 _04435_ net1169 vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__o211a_1
XANTENNA__16222__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11363_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] team_01_WB.instance_to_wrap.cpu.f0.i\[17\]
+ _07690_ vssd1 vssd1 vccd1 vccd1 _07692_ sky130_fd_sc_hd__and3_1
X_13102_ net56 net55 net58 net57 vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__or4_1
X_10314_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[18\] net945
+ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__and3_1
X_14082_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[76\] _04235_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[76\]
+ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__a22o_1
X_11294_ _04714_ _07627_ _04734_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1
+ vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17910_ net1602 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
X_13033_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[53\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[61\]
+ net855 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10245_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[9\] net777 net755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__a22o_1
XANTENNA__12290__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1100 net1105 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__buf_2
XFILLER_0_119_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16372__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1111 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[22\] vssd1 vssd1 vccd1 vccd1
+ net1111 sky130_fd_sc_hd__buf_2
X_10176_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[10\] net779 _06514_
+ _06515_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__a211o_1
X_17841_ clknet_leaf_77_wb_clk_i net2576 _01781_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[111\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1122 net1126 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09751__A2 _04636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14088__A1 _04348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1133 net1135 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__buf_2
Xfanout1144 net1145 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__clkbuf_2
Xfanout1155 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1 vccd1
+ net1155 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1166 net1167 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__buf_2
X_17772_ clknet_leaf_68_wb_clk_i net1668 _01712_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10104__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14984_ net1289 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__inv_2
Xfanout1177 net1204 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__clkbuf_2
Xfanout190 net192 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_2
Xfanout1188 net1194 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1199 net1202 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__buf_4
XANTENNA__10649__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13935_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__and2b_2
X_16723_ clknet_leaf_135_wb_clk_i _02410_ _00706_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16654_ clknet_leaf_8_wb_clk_i _02341_ _00637_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13866_ net1164 net1059 net3283 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[27\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_53_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08509__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15605_ net1219 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12817_ net1650 net640 net607 _03640_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a22o_1
X_16585_ clknet_leaf_14_wb_clk_i _02272_ _00568_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_13797_ _04175_ _04178_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15536_ net1270 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__inv_2
X_12748_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] net1054 net363 _03592_
+ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15467_ net1298 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__inv_2
XANTENNA__12465__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08490__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12679_ net2055 net281 net390 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__mux2_1
XANTENNA__14246__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17206_ clknet_leaf_141_wb_clk_i _02893_ _01189_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14418_ net1365 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15398_ net1325 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17137_ clknet_leaf_18_wb_clk_i _02824_ _01120_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_113_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14349_ net1375 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__inv_2
Xhold605 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire591 _04880_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__clkbuf_1
Xhold616 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold627 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17068_ clknet_leaf_133_wb_clk_i _02755_ _01051_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09990__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11809__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08910_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[2\] net672 _05229_ _05239_
+ _05246_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_100_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15077__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16019_ net1377 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09890_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[5\] net946 vssd1
+ vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08841_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[1\] net695 _05156_ _05157_
+ _05170_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09506__C net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1305 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1316 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2932 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16865__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1327 _02150_ vssd1 vssd1 vccd1 vccd1 net2943 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15805__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08772_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] net730 _05111_ net1105 vssd1
+ vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1338 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1349 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout344_A _04748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1086_A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09324_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[24\] net687 net673 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__a22o_1
XANTENNA__15540__A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10812__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09255_ net598 _05591_ _05593_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__o21a_1
XANTENNA__12375__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout511_A _05963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1253_A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08206_ net2867 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[67\] net1051 vssd1 vssd1
+ vccd1 vccd1 _03481_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_90_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09186_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[16\] net685 _05523_
+ _05524_ _05525_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12565__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13995__A _04152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08137_ _04467_ team_01_WB.instance_to_wrap.cpu.f0.num\[28\] team_01_WB.instance_to_wrap.cpu.f0.num\[21\]
+ _04473_ _04596_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10576__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_83_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09981__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ _04514_ _04532_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout880_A _04810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17640__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11719__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12868__A2 _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[0\] net975 vssd1
+ vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__and3_1
XANTENNA__09733__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17790__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ net2547 net253 net472 vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13720_ _04107_ _04129_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[11\]
+ sky130_fd_sc_hd__nor2_1
X_10932_ _05338_ _06563_ vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18075__1575 vssd1 vssd1 vccd1 vccd1 _18075__1575/HI net1575 sky130_fd_sc_hd__conb_1
XFILLER_0_54_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08329__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17020__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13651_ _03877_ _03879_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__xnor2_1
X_10863_ _06980_ _07132_ _07202_ _06920_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_116_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12602_ net2290 net235 net395 vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__mux2_1
X_16370_ clknet_leaf_62_wb_clk_i _02124_ _00353_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[93\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13889__B _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13582_ net723 _07541_ net1068 vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__o21a_1
X_10794_ _06963_ _07122_ _07133_ _07054_ _07131_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08990__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15321_ net1259 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12533_ net3178 net245 net403 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12285__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10594__A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17170__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18040_ net1540 vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__buf_2
XFILLER_0_87_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15252_ net1268 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12464_ net2849 net276 net413 vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__mux2_1
XANTENNA__16738__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14203_ net1677 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11415_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] _07705_ vssd1 vssd1 vccd1 vccd1
+ _07731_ sky130_fd_sc_hd__or2_1
XANTENNA__11202__B _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15183_ net1214 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__inv_2
XANTENNA__10567__A0 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12395_ net3146 net213 net419 vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08999__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14134_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[31\] _04243_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[119\]
+ _04418_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__a221o_1
XANTENNA__09972__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11346_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] team_01_WB.instance_to_wrap.cpu.f0.i\[4\]
+ _07674_ vssd1 vssd1 vccd1 vccd1 _07675_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_91_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14065_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[19\] _04259_ _04349_ _04351_
+ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__a2111o_1
XANTENNA__16888__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10319__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ _05595_ net332 _07354_ net337 net370 vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13016_ net2262 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[78\] net852 vssd1 vssd1
+ vccd1 vccd1 _02109_ sky130_fd_sc_hd__mux2_1
X_10228_ _06566_ _06567_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__nand2_1
XANTENNA__11531__A2 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_135_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17824_ clknet_leaf_75_wb_clk_i net2518 _01764_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10159_ _06497_ _06498_ net341 vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__a21oi_1
Xhold2 team_01_WB.instance_to_wrap.cpu.RU0.state\[1\] vssd1 vssd1 vccd1 vccd1 net1618
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17755_ clknet_leaf_71_wb_clk_i _03431_ _01695_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14967_ net1195 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16706_ clknet_leaf_35_wb_clk_i _02393_ _00689_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10098__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13918_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\] _04212_ net572 vssd1
+ vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_102_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14898_ net1233 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17686_ clknet_leaf_94_wb_clk_i _03370_ _01627_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_134_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16637_ clknet_leaf_50_wb_clk_i _02324_ _00620_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09061__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13849_ net1166 net1060 net2152 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[10\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__16268__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16568_ clknet_leaf_25_wb_clk_i _02255_ _00551_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_80_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12795__A1 _07207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13992__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12195__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15519_ net1260 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16499_ clknet_leaf_105_wb_clk_i _02253_ _00482_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09040_ net1155 net619 net593 vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_2_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17663__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold402 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[20\] vssd1 vssd1 vccd1 vccd1
+ net2018 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold413 net123 vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10022__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold424 team_01_WB.instance_to_wrap.cpu.f0.i\[7\] vssd1 vssd1 vccd1 vccd1 net2040
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13441__A_N _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold468 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ net378 _05264_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold479 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout904 net905 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__buf_4
XFILLER_0_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12224__A _07784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout915 net916 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09715__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout926 net928 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_8
X_09873_ _06198_ _06210_ _06211_ _06212_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__or4_1
Xfanout937 _04759_ vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__buf_4
Xfanout948 net950 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__buf_4
XANTENNA_fanout294_A _07926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 _04650_ vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__buf_4
X_08824_ net1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[1\] net887 vssd1
+ vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__and3_1
Xhold1102 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[94\] vssd1 vssd1 vccd1 vccd1
+ net2718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2729 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1001_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2762 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09533__A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08755_ net1088 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[4\] net920 vssd1
+ vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__and3_1
Xhold1157 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2773 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout461_A _07955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1168 team_01_WB.instance_to_wrap.cpu.f0.num\[9\] vssd1 vssd1 vccd1 vccd1 net2784
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1179 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2795 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10089__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_130_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08686_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[7\] net882 vssd1
+ vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout726_A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1370_A net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09307_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[22\] net675 _05621_
+ _05631_ _05639_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12786__A1 _07188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13983__B1 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10797__A0 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11303__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09238_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[21\] net697 net696 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[21\]
+ _05577_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_40_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08315__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11022__B net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[16\] net653 _05506_
+ _05507_ _05508_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10549__A0 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09403__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ _06963_ _07054_ _07324_ net555 vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10013__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ net3035 net285 net450 vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11131_ _06399_ _06401_ vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_129_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11062_ _07394_ _07398_ _07400_ _07401_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10013_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[1\] net781 net763 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15870_ net1350 vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_34_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08985__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ net1207 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__inv_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10589__A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16410__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17536__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17540_ clknet_leaf_54_wb_clk_i _03227_ _01523_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14752_ net1315 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11964_ net2520 net215 net473 vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11277__B2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13703_ _04104_ _04119_ _04122_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[7\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__08142__B2 _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10915_ net375 net374 _06738_ _06158_ net539 net546 vssd1 vssd1 vccd1 vccd1 _07255_
+ sky130_fd_sc_hd__mux4_1
X_17471_ clknet_leaf_24_wb_clk_i _03158_ _01454_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14683_ net1344 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11895_ net2448 net220 net479 vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__mux2_1
XANTENNA__08693__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11912__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16422_ clknet_leaf_106_wb_clk_i _02176_ _00405_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13634_ net724 _07290_ team_01_WB.instance_to_wrap.cpu.IM0.pc_enable vssd1 vssd1
+ vccd1 vccd1 _04072_ sky130_fd_sc_hd__o21a_1
X_10846_ net529 _06921_ _06972_ _06978_ _07185_ vssd1 vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_6_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16560__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17686__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16353_ clknet_leaf_57_wb_clk_i _02107_ _00336_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[76\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_15_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13412__B _05224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13565_ net722 _07135_ net1066 vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__o21a_1
X_10777_ net509 net508 net507 net505 net548 net538 vssd1 vssd1 vccd1 vccd1 _07117_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15304_ net1283 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12516_ net1828 net294 net410 vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16284_ clknet_leaf_94_wb_clk_i _02038_ _00267_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13496_ net186 _03955_ _03956_ net726 vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18023_ net1523 vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__buf_2
XFILLER_0_129_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15235_ net1187 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__inv_2
X_12447_ net2822 _07912_ net417 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15166_ net1275 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__inv_2
X_12378_ net2554 net228 net425 vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__mux2_1
XANTENNA__08522__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14117_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[110\] _04264_ _04400_ _04402_
+ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11329_ _04547_ _07653_ _07662_ net1162 vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__a2bb2o_1
X_15097_ net1259 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__inv_2
XANTENNA__10490__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17066__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14048_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[67\] _04233_ _04260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[59\]
+ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09056__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11504__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08895__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17807_ clknet_leaf_61_wb_clk_i _03483_ _01747_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[77\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_136_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15999_ net1405 vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11268__A1 _06915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08540_ _04871_ _04872_ _04878_ _04879_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__nor4_1
XANTENNA__11268__B2 _06912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17738_ clknet_leaf_84_wb_clk_i _03414_ _01678_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13662__C1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09330__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16903__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08471_ net1086 net879 vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17669_ clknet_leaf_117_wb_clk_i _03354_ _01610_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15090__A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11822__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12768__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11123__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17921__1609 vssd1 vssd1 vccd1 vccd1 net1609 _17921__1609/LO sky130_fd_sc_hd__conb_1
XFILLER_0_17_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09023_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[9\] net690 _05342_ _05347_
+ _05362_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_86_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12653__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout307_A _07935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1049_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 _02021_ vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold221 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[5\] vssd1 vssd1 vccd1 vccd1 net1837
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09936__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17409__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08432__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold232 team_01_WB.instance_to_wrap.a1.ADR_I\[21\] vssd1 vssd1 vccd1 vccd1 net1848
+ sky130_fd_sc_hd__dlygate4sd3_1
X_18074__1574 vssd1 vssd1 vccd1 vccd1 _18074__1574/HI net1574 sky130_fd_sc_hd__conb_1
XFILLER_0_41_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12940__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold243 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[27\] vssd1 vssd1 vccd1 vccd1 net1859
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold254 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1
+ net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 team_01_WB.instance_to_wrap.cpu.c0.count\[10\] vssd1 vssd1 vccd1 vccd1 net1881
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold276 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1216_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold287 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout701 _04760_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_4
X_09925_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[4\] net791 _06262_ _06263_
+ _06264_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14142__B1 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold298 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout712 net713 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__clkbuf_4
Xfanout723 net724 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__clkbuf_4
Xfanout734 _04688_ vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__buf_4
XANTENNA_fanout676_A _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 _04684_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_8
Xfanout756 _04675_ vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__buf_6
XANTENNA__16433__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17559__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout767 _04673_ vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__clkbuf_8
X_09856_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[12\] net796 net777 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__a22o_1
Xfanout778 _04666_ vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__buf_8
Xfanout789 net790 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_8
X_08807_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[0\] net879 vssd1
+ vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__and3_1
Xclkbuf_4_8__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09787_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\] net765 vssd1 vssd1
+ vccd1 vccd1 _06127_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout843_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ net1088 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[4\] net881 vssd1
+ vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10202__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13653__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09321__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08669_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[7\] net893 vssd1
+ vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_137_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10700_ net534 _06955_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11680_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[15\] net717 vssd1 vssd1 vccd1
+ vccd1 _07881_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12759__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10631_ net515 net503 vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08326__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17933__1435 vssd1 vssd1 vccd1 vccd1 _17933__1435/HI net1435 sky130_fd_sc_hd__conb_1
XFILLER_0_14_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10234__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ team_01_WB.instance_to_wrap.cpu.f0.i\[11\] _07677_ vssd1 vssd1 vccd1 vccd1
+ _03823_ sky130_fd_sc_hd__or2_1
X_10562_ _06900_ _06901_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__or2_2
XFILLER_0_24_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12301_ net2896 net201 net431 vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13281_ _07650_ _03767_ _03769_ net825 net1631 vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__o32a_1
XANTENNA__12563__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10493_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[31\] net959 vssd1
+ vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__and3b_1
XFILLER_0_121_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15020_ net1180 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12232_ net2486 net209 net441 vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__mux2_1
XANTENNA__08342__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12931__A1 _05453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12163_ net2614 net248 net448 vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__mux2_1
XANTENNA__10942__A0 _06636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ _07452_ _07453_ net541 vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__mux2_1
XANTENNA__14133__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16971_ clknet_leaf_0_wb_clk_i _02658_ _00954_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12094_ net2866 net221 net457 vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11907__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11045_ _05189_ _07011_ _06366_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15922_ net1331 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09173__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15853_ net1363 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09604__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14804_ net1291 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__inv_2
X_12996_ net2817 net2599 net859 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15784_ net1307 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17523_ clknet_leaf_135_wb_clk_i _03210_ _01506_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11947_ net1895 net254 net476 vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14735_ net1321 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11642__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17454_ clknet_leaf_5_wb_clk_i _03141_ _01437_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14666_ net1376 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11878_ net2058 net257 net484 vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08517__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16405_ clknet_leaf_79_wb_clk_i _02159_ _00388_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13617_ net723 _07207_ net1068 vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__o21a_1
X_10829_ _07064_ _07099_ _07167_ _07168_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14597_ net1403 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__inv_2
X_17385_ clknet_leaf_9_wb_clk_i _03072_ _01368_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16306__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16336_ clknet_leaf_71_wb_clk_i _02090_ _00319_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_13548_ net722 _07154_ net1066 vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16267_ clknet_leaf_104_wb_clk_i net1791 _00255_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10782__A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13479_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _05679_ vssd1 vssd1
+ vccd1 vccd1 _03940_ sky130_fd_sc_hd__xor2_1
XANTENNA__12473__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18006_ net1506 vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_hd__buf_2
X_15218_ net1232 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09379__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09918__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16198_ clknet_leaf_114_wb_clk_i _01958_ _00186_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15149_ net1215 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10933__A0 _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17701__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14124__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07971_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1 _04469_
+ sky130_fd_sc_hd__inv_2
XANTENNA__11817__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09710_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[21\] net794 _06038_ _06039_
+ _06040_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__a2111o_1
XANTENNA__15085__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[23\] net811 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17851__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09572_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[25\] net970
+ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08523_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[18\] net900
+ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__and3_1
XANTENNA__12648__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08657__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11110__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout257_A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13650__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08454_ net1024 net894 vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__and2_1
XANTENNA__10464__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11661__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08385_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout424_A _07966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1166_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17231__CLK clknet_leaf_143_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12383__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09006_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[9\] net898 vssd1
+ vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__and3_1
XANTENNA__13166__B2 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09909__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08042__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14115__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16949__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout520 net521 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_2
Xfanout531 net532 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_4
Xfanout542 _05189_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__buf_2
X_09908_ net770 _06240_ _06244_ _06247_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__or4_2
Xfanout553 _05115_ vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__buf_2
Xfanout564 net566 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout575 _07792_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout586 _04517_ vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_4
X_09839_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[13\] net815 net739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__a22o_1
Xfanout597 _04840_ vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12850_ net3094 net233 net380 vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ net2891 net203 net491 vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12558__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12781_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] net1056 net365 _03615_
+ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ net1383 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11732_ net718 _07507_ net613 vssd1 vssd1 vccd1 vccd1 _07923_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10455__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14451_ net1374 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__inv_2
X_11663_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] _07812_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\]
+ vssd1 vssd1 vccd1 vccd1 _07868_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_94_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\]
+ net596 vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__and3_1
XANTENNA__10207__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10614_ net547 _06366_ vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__nor2_1
X_17170_ clknet_leaf_129_wb_clk_i _02857_ _01153_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14382_ net1304 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09073__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11594_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _07809_ vssd1 vssd1
+ vccd1 vccd1 _07811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16121_ clknet_leaf_100_wb_clk_i _01896_ _00109_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13333_ team_01_WB.instance_to_wrap.cpu.f0.i\[15\] _07682_ net827 vssd1 vssd1 vccd1
+ vccd1 _03810_ sky130_fd_sc_hd__o21a_1
XANTENNA__12293__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10545_ _06883_ _06884_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08820__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17724__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09168__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16052_ clknet_leaf_89_wb_clk_i _01845_ _00040_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13264_ net586 _03750_ _03755_ net565 _04466_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_121_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10476_ _05931_ _05933_ _05963_ _05964_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__a22o_1
XANTENNA__08072__A team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12904__A1 _05591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15003_ net1180 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__inv_2
XANTENNA__11707__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ net2483 net279 net443 vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08033__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10915__A0 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13195_ net14 net835 net628 net2160 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14106__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ net2370 net253 net453 vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09781__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17874__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11637__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16954_ clknet_leaf_60_wb_clk_i _02641_ _00937_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12077_ net2999 net255 net460 vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15905_ net1337 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11028_ _07366_ _07367_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16885_ clknet_leaf_123_wb_clk_i _02572_ _00868_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_17920__1608 vssd1 vssd1 vccd1 vccd1 net1608 _17920__1608/LO sky130_fd_sc_hd__conb_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17104__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11891__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15836_ net1370 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13093__A0 _03716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09631__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12979_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[107\] net3057 net865 vssd1 vssd1
+ vccd1 vccd1 _02146_ sky130_fd_sc_hd__mux2_1
XANTENNA__12468__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15767_ net1346 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__inv_2
XANTENNA__13632__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18073__1573 vssd1 vssd1 vccd1 vccd1 _18073__1573/HI net1573 sky130_fd_sc_hd__conb_1
XFILLER_0_38_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17506_ clknet_leaf_34_wb_clk_i _03193_ _01489_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14718_ net1315 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__inv_2
XANTENNA__11643__A1 _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15698_ net1235 vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__inv_2
XANTENNA__17254__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17437_ clknet_leaf_20_wb_clk_i _03124_ _01420_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14649_ net1174 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_16 _06737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_27 _07873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ net2575 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[103\] net1047 vssd1 vssd1
+ vccd1 vccd1 _03517_ sky130_fd_sc_hd__mux2_1
XANTENNA_49 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17368_ clknet_leaf_28_wb_clk_i _03055_ _01351_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16319_ clknet_leaf_66_wb_clk_i _02073_ _00302_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08811__A2 _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17299_ clknet_leaf_129_wb_clk_i _02986_ _01282_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
XFILLER_0_3_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09509__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XANTENNA__15808__A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
XANTENNA__13182__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_112_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
XANTENNA__09772__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput178 net178 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XANTENNA__08710__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10382__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17932__1434 vssd1 vssd1 vccd1 vccd1 _17932__1434/HI net1434 sky130_fd_sc_hd__conb_1
XANTENNA_fanout374_A _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09624_ _05682_ _05734_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09541__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13084__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09555_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[28\] net792 net770 _05883_
+ _05894_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_37_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12378__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1283_A net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13623__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ net712 _04838_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__or2_2
XANTENNA__11634__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12831__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[30\] net677 net649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08437_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[23\] net915 vssd1
+ vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16621__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_A _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08368_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\] _04623_ _04626_ vssd1 vssd1
+ vccd1 vccd1 _04708_ sky130_fd_sc_hd__nor3_2
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08299_ net989 net969 vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10330_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] net765 net621 vssd1
+ vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11030__B net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10261_ _06590_ _06593_ _06566_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__a21boi_2
XANTENNA__12841__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12000_ net3007 net276 net469 vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10192_ _06530_ _06531_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__or2_1
Xfanout1304 net1305 vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__buf_4
Xfanout1315 net1317 vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__buf_4
XANTENNA__17127__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1326 net1329 vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__buf_2
Xfanout1337 net1340 vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__clkbuf_4
Xfanout1348 net1349 vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__buf_4
Xfanout350 _03742_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_2
Xfanout361 _03653_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_2
Xfanout1359 net1414 vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__buf_2
Xfanout372 _06738_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_2
X_13951_ _04225_ _04242_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__nor2_4
Xfanout383 _03570_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_6
XANTENNA__10125__B2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08869__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout394 _03568_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12902_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[22\] net1031 vssd1 vssd1 vccd1
+ vccd1 _03677_ sky130_fd_sc_hd__or2_1
X_13882_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[4\]
+ _04188_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__and3_2
X_16670_ clknet_leaf_48_wb_clk_i _02357_ _00653_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16151__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17277__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08993__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15621_ net1208 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12833_ net575 _07794_ _07945_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__and3_1
XANTENNA__12288__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09818__A1 _06157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10428__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15552_ net1243 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__inv_2
X_12764_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[21\] _07621_ net1025 vssd1 vssd1
+ vccd1 vccd1 _03604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14503_ net1329 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__inv_2
XANTENNA__10979__A3 _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11715_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[8\] _07290_ net719 vssd1 vssd1
+ vccd1 vccd1 _07909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15483_ net1181 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__inv_2
X_12695_ net2561 net276 net385 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__mux2_1
XANTENNA__11920__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17222_ clknet_leaf_38_wb_clk_i _02909_ _01205_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14434_ net1396 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__inv_2
X_11646_ _07852_ _07854_ net611 vssd1 vssd1 vccd1 vccd1 _07855_ sky130_fd_sc_hd__mux2_4
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17153_ clknet_leaf_41_wb_clk_i _02840_ _01136_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
X_14365_ net1353 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput36 gpio_in[18] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
X_11577_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\]
+ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__and2_2
XFILLER_0_13_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput47 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__buf_1
X_13316_ net565 _07708_ _03796_ net829 vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__a31o_1
X_16104_ clknet_leaf_91_wb_clk_i _01879_ _00092_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput58 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
X_17084_ clknet_leaf_37_wb_clk_i _02771_ _01067_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput69 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
X_10528_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[31\] net683 net668 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold809 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[115\] vssd1 vssd1 vccd1 vccd1
+ net2425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14296_ net1355 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16035_ clknet_leaf_103_wb_clk_i _01829_ _00029_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13247_ net2000 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1
+ vccd1 vccd1 _01903_ sky130_fd_sc_hd__a22o_1
X_10459_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[26\] net813 net776 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09754__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13550__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09626__A _05963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ net107 net844 net631 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__a21o_1
XANTENNA__08530__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12129_ net2433 net215 net451 vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17986_ net1486 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_40_1450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1509 team_01_WB.instance_to_wrap.a1.ADR_I\[6\] vssd1 vssd1 vccd1 vccd1 net3125
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16937_ clknet_leaf_10_wb_clk_i _02624_ _00920_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09064__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16868_ clknet_leaf_54_wb_clk_i _02555_ _00851_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15819_ net1314 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__inv_2
XANTENNA__12198__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16799_ clknet_leaf_26_wb_clk_i _02486_ _00782_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16644__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09340_ net601 _05679_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__or2_1
XANTENNA__11616__A1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12813__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10300__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09271_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[20\] net663 net659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11830__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ net3064 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[51\] net1051 vssd1 vssd1
+ vccd1 vccd1 _03465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_80_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08705__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14030__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08153_ net1750 net826 _00020_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08084_ _04528_ _04532_ _04527_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12661__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1031_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1129_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13541__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_A _07944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout589_A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[8\] net879 vssd1
+ vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__and3_1
XANTENNA__14097__A2 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16174__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout756_A _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09607_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[24\] net944 vssd1
+ vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09702__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout923_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09538_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[28\] net944
+ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09276__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11025__B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09469_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[30\] net878
+ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__and3_1
XANTENNA__11083__A2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12836__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11500_ net1846 net876 _07758_ _07777_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__o22a_1
XFILLER_0_65_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12480_ net3262 net303 net412 vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09028__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14021__A2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11431_ _07680_ _07701_ _07740_ net327 vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_134_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08334__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10043__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14055__C _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14150_ _04422_ _04431_ _04433_ _04434_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11362_ team_01_WB.instance_to_wrap.cpu.f0.i\[17\] _07690_ vssd1 vssd1 vccd1 vccd1
+ _07691_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13101_ net47 net49 net48 net46 vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__or4b_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10313_ _06650_ _06651_ _06652_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__or3_1
X_14081_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[124\] _04263_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[108\]
+ _04368_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__a221o_1
XANTENNA__12571__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11293_ _07627_ _07629_ _07632_ vssd1 vssd1 vccd1 vccd1 _07633_ sky130_fd_sc_hd__a21boi_1
X_13032_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[54\] net2359 net853 vssd1 vssd1
+ vccd1 vccd1 _02093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10244_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[9\] net823 net787 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__a22o_1
XANTENNA__08988__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18072__1572 vssd1 vssd1 vccd1 vccd1 _18072__1572/HI net1572 sky130_fd_sc_hd__conb_1
XANTENNA__16517__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11695__B net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09446__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input52_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1101 net1104 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__buf_2
X_17840_ clknet_leaf_75_wb_clk_i _03516_ _01780_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1112 net1113 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_125_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10175_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[10\] net785 net739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1123 net1126 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14088__A2 _04375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1134 net1135 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1145 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1 vccd1 vccd1
+ net1145 sky130_fd_sc_hd__clkbuf_2
Xfanout1156 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[6\] vssd1 vssd1 vccd1 vccd1
+ net1156 sky130_fd_sc_hd__buf_2
X_17771_ clknet_leaf_70_wb_clk_i _03447_ _01711_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[41\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1167 net3185 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__clkbuf_2
X_14983_ net1301 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__inv_2
XANTENNA__13296__B1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1178 net1182 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__buf_4
XANTENNA__11915__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16667__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 net192 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__buf_2
Xfanout1189 net1194 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__buf_2
X_16722_ clknet_leaf_131_wb_clk_i _02409_ _00705_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13934_ _04224_ _04225_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__nor2_4
XFILLER_0_96_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09181__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16653_ clknet_leaf_140_wb_clk_i _02340_ _00636_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13865_ net1163 net1059 net2233 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[26\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_44_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15604_ net1268 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12816_ net366 _03638_ _03639_ net1057 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__a32o_1
XFILLER_0_134_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16584_ clknet_leaf_24_wb_clk_i _02271_ _00567_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13796_ _04177_ _04174_ _01836_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__mux2_1
XANTENNA__09267__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15535_ net1216 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[26\] _07588_ net1026 vssd1 vssd1
+ vccd1 vccd1 _03592_ sky130_fd_sc_hd__mux2_1
XANTENNA__11650__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10282__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12678_ net2941 net302 net390 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__mux2_1
X_15466_ net1278 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__inv_2
XANTENNA__14012__A2 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08525__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17205_ clknet_leaf_126_wb_clk_i _02892_ _01188_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12023__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14417_ net1360 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__inv_2
X_11629_ _07819_ _07840_ vssd1 vssd1 vccd1 vccd1 _07841_ sky130_fd_sc_hd__nor2_1
X_17931__1433 vssd1 vssd1 vccd1 vccd1 _17931__1433/HI net1433 sky130_fd_sc_hd__conb_1
XANTENNA__13840__A_N net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15397_ net1205 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10493__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17136_ clknet_leaf_127_wb_clk_i _02823_ _01119_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14348_ net1357 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09059__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold606 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10585__A1 _06882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire581 _06705_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_2
Xhold617 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 net2233
+ sky130_fd_sc_hd__dlygate4sd3_1
Xwire592 _04877_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold628 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[17\] vssd1 vssd1 vccd1 vccd1
+ net2244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[15\] vssd1 vssd1 vccd1 vccd1
+ net2255 sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ net1367 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__inv_2
X_17067_ clknet_leaf_5_wb_clk_i _02754_ _01050_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12481__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16197__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13523__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08898__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16018_ net1357 vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11534__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08840_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[1\] net664 _05159_ _05173_
+ _05174_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14079__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1306 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[41\] vssd1 vssd1 vccd1 vccd1
+ net2922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1317 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2933 sky130_fd_sc_hd__dlygate4sd3_1
X_08771_ _04708_ net726 net720 _04838_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__or4_2
Xhold1328 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2944 sky130_fd_sc_hd__dlygate4sd3_1
X_17969_ net1469 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
XANTENNA__13287__B1 _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1339 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17592__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08702__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10030__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09258__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09323_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[24\] net697 net677 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__a22o_1
XANTENNA__12656__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout337_A _06911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09254_ net598 _05591_ _05593_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout1079_A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14003__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08205_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[76\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[68\]
+ net1041 vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09185_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[16\] net913
+ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__and3_1
XANTENNA__13211__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout504_A _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1246_A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] _04494_ team_01_WB.instance_to_wrap.cpu.f0.num\[0\]
+ _04489_ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10576__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09430__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ _04528_ _04539_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__nor2_1
XANTENNA__12391__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1413_A net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13514__A1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14900__A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13278__B1 _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[8\] net885 vssd1
+ vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_51_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ net2645 net227 net472 vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10931_ _05338_ _06563_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08329__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10862_ net503 _07105_ net376 vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13650_ net983 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] _04083_ _04084_
+ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09249__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12601_ net3118 net239 net395 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__mux2_1
X_13581_ net188 _04025_ _04026_ net729 vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__a211o_1
X_10793_ net528 _07132_ _07119_ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12566__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13889__C _04195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17315__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15320_ net1176 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__inv_2
X_12532_ net3205 net201 net403 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08345__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10594__B _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15251_ net1281 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12463_ net2049 net210 net414 vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__mux2_1
XANTENNA__13202__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10016__B1 _04687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14202_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\] vssd1 vssd1 vccd1
+ vccd1 _02285_ sky130_fd_sc_hd__clkbuf_1
X_11414_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] _07691_ vssd1 vssd1 vccd1 vccd1
+ _07730_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15182_ net1284 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12394_ net2776 net217 net419 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__mux2_1
XANTENNA__11202__C _07531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09421__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10567__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[47\] _04246_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[111\]
+ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11345_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] _07673_ vssd1 vssd1 vccd1 vccd1
+ _07674_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09709__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14064_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[11\] _04253_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[115\]
+ _04352_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__a221o_1
XANTENNA__09176__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ _06919_ _07354_ vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__nor2_1
XANTENNA__09607__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ net2498 net2435 net861 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__mux2_1
XANTENNA__08511__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10227_ _06562_ _06565_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__or2_1
X_17823_ clknet_leaf_61_wb_clk_i _03499_ _01763_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[93\]
+ sky130_fd_sc_hd__dfstp_1
X_10158_ net378 _05379_ net377 vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__a21o_1
Xhold3 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[19\] vssd1 vssd1 vccd1 vccd1 net1619
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17754_ clknet_leaf_76_wb_clk_i net2008 _01694_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14966_ net1201 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__inv_2
X_10089_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[7\] net785 net782 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_106_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16705_ clknet_leaf_42_wb_clk_i _02392_ _00688_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13917_ _04212_ net572 _04211_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_102_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17685_ clknet_leaf_94_wb_clk_i _03369_ _01626_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_102_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14897_ net1289 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
X_16636_ clknet_leaf_37_wb_clk_i _02323_ _00619_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13848_ net1166 net1060 net1672 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[9\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12476__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16567_ clknet_leaf_108_wb_clk_i net833 _00550_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.ihit
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_58_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13779_ net1170 _04163_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14257__A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15518_ net1252 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16498_ clknet_leaf_104_wb_clk_i _02252_ _00481_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17808__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15449_ net1258 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__inv_2
XANTENNA__10007__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11755__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09412__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[3\] vssd1 vssd1 vccd1 vccd1
+ net2019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 _01989_ vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
X_17119_ clknet_leaf_8_wb_clk_i _02806_ _01102_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08620__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold425 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
X_18099_ net1588 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_0_64_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold447 team_01_WB.instance_to_wrap.a1.ADR_I\[8\] vssd1 vssd1 vccd1 vccd1 net2063
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09086__A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold458 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold469 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ _06280_ vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_74_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12224__B _07789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08421__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout905 _04785_ vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout916 net918 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_8
Xfanout927 net928 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__buf_4
X_09872_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[12\] net798 net758 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__a22o_1
Xfanout938 net940 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__buf_6
Xfanout949 net950 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_2
X_08823_ net1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[1\] net927 vssd1
+ vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__and3_1
Xhold1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2719 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16982__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1114 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2730 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_7__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xhold1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2752 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ net1008 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[4\] net901 vssd1
+ vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__and3_1
Xhold1147 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2774 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1169 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2785 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09479__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08685_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[7\] net910 vssd1
+ vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__and3_1
XANTENNA__16212__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17338__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12386__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18071__1571 vssd1 vssd1 vccd1 vccd1 _18071__1571/HI net1571 sky130_fd_sc_hd__conb_1
XANTENNA_fanout621_A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1363_A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09306_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[22\] net655 _05628_
+ _05642_ _05643_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_64_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout719_A _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16362__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09651__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17488__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10797__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09237_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[21\] net694 net662 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_131_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11303__B _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09939__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09168_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[16\] net885 vssd1
+ vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10549__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout990_A _04491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08119_ _04483_ team_01_WB.instance_to_wrap.cpu.f0.num\[10\] team_01_WB.instance_to_wrap.cpu.f0.num\[5\]
+ _04488_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_62_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09099_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[13\] net894 vssd1
+ vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__and3_1
XANTENNA__08611__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11130_ _06920_ _07216_ _07228_ _06928_ net330 vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold970 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[99\] vssd1 vssd1 vccd1 vccd1
+ net2586 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold981 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14160__A1 _04195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold992 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[74\] vssd1 vssd1 vccd1 vccd1
+ net2608 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ _05042_ _06438_ _07381_ _07399_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_25_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10012_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[1\] net817 net797 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ net1239 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17930__1432 vssd1 vssd1 vccd1 vccd1 _17930__1432/HI net1432 sky130_fd_sc_hd__conb_1
XANTENNA__10589__B _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1670 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 net3286
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14751_ net1315 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__inv_2
XANTENNA__11277__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09162__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11963_ net2417 net216 net471 vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13671__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13702_ team_01_WB.instance_to_wrap.cpu.c0.count\[7\] _04103_ vssd1 vssd1 vccd1 vccd1
+ _04122_ sky130_fd_sc_hd__or2_1
X_17470_ clknet_leaf_45_wb_clk_i _03157_ _01453_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10914_ net342 net341 _06526_ net340 net551 net542 vssd1 vssd1 vccd1 vccd1 _07254_
+ sky130_fd_sc_hd__mux4_1
X_14682_ net1361 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__inv_2
X_11894_ net3258 net223 net479 vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16421_ clknet_leaf_106_wb_clk_i _02175_ _00404_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10845_ _06921_ _06965_ vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__or2_2
XFILLER_0_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13633_ net187 _04069_ _04070_ net728 vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12296__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10237__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16352_ clknet_leaf_74_wb_clk_i _02106_ _00335_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11434__C1 _07699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13564_ net185 _04011_ _04012_ net726 vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__a211o_1
X_10776_ _06641_ _06675_ _07114_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__nand3_1
XANTENNA__08075__A team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10788__A1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09642__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15303_ net1327 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__inv_2
X_12515_ net2150 net301 net410 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16283_ clknet_leaf_56_wb_clk_i _02037_ _00266_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13495_ net198 net194 _07822_ net644 vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_114_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16855__CLK clknet_leaf_137_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18022_ net1522 vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__buf_2
XFILLER_0_136_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13726__A1 team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12446_ net3020 net286 net417 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__mux2_1
X_15234_ net1266 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12377_ net2375 net289 net425 vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15165_ net1251 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14116_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[62\] _04258_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[126\]
+ _04401_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__a221o_1
X_11328_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] _07659_ vssd1 vssd1 vccd1
+ vccd1 _07662_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_26_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15096_ net1183 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__inv_2
X_14047_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[11\] _04226_ _04244_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[99\]
+ _04335_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__a221o_1
X_11259_ _06935_ _07281_ _07597_ _07598_ vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_108_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09634__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16235__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17806_ clknet_leaf_57_wb_clk_i _03482_ _01746_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[76\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15998_ net1395 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17737_ clknet_leaf_81_wb_clk_i net1749 _01677_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14949_ net1205 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10476__B1 _05963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08470_ net1109 net1114 net1112 net1106 vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_89_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17668_ clknet_leaf_117_wb_clk_i _03353_ _01609_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16385__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16619_ clknet_leaf_5_wb_clk_i _02306_ _00602_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17599_ clknet_leaf_70_wb_clk_i _03286_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12768__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09022_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[9\] net890 vssd1
+ vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08713__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09397__A1 _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13193__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold200 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[7\] vssd1 vssd1 vccd1 vccd1
+ net1816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout202_A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold222 _01971_ vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08432__B net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold233 _02019_ vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _01993_ vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12940__A2 _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold255 net117 vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold266 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[122\] vssd1 vssd1 vccd1 vccd1
+ net1904 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[4\] net944 vssd1
+ vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__and3_1
Xfanout702 _04758_ vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_8
Xhold299 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout713 _04728_ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout724 _04721_ vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1209_A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout735 _04687_ vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__clkbuf_8
Xfanout746 _04682_ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__buf_6
X_09855_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[12\] net780 net754 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__a22o_1
Xfanout757 _04675_ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 _04672_ vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10703__A1 _07042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout779 net781 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_8
X_18089__1586 vssd1 vssd1 vccd1 vccd1 _18089__1586/HI net1586 sky130_fd_sc_hd__conb_1
XANTENNA__17160__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[0\] net885 vssd1
+ vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09786_ net770 _06119_ _06122_ _06125_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__or4_1
XFILLER_0_55_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08737_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[4\] net920 vssd1
+ vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout836_A _03737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08668_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[7\] net889 vssd1
+ vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09872__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[15\] net671 _04937_ _04938_
+ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__a211o_1
XANTENNA__13005__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10219__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ net533 net503 vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10561_ _04736_ _04738_ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12844__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11431__A2 _07701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12300_ net2484 net207 net431 vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13280_ _03754_ _03768_ _04621_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10492_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[31\] net952
+ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12231_ net3078 net247 net441 vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__mux2_1
XANTENNA__13184__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08342__B net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12931__A2 _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ net2954 net213 net448 vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09157__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10942__A1 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11113_ _06947_ _06951_ vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__nor2_1
XANTENNA__16258__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12093_ net3271 net223 net455 vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__mux2_1
X_16970_ clknet_leaf_11_wb_clk_i _02657_ _00953_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15921_ net1339 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__inv_2
X_11044_ _07382_ _07383_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__nand2b_1
XANTENNA__11498__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08363__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15852_ net1364 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__inv_2
XANTENNA__10170__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14803_ net1233 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__inv_2
XANTENNA__12447__A1 _07912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15783_ net1306 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__inv_2
XANTENNA__13644__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12995_ net2383 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[99\] net865 vssd1 vssd1
+ vccd1 vccd1 _02130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11923__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17522_ clknet_leaf_130_wb_clk_i _03209_ _01505_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14734_ net1318 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11946_ net2265 net228 net475 vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09863__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17453_ clknet_leaf_140_wb_clk_i _03140_ _01436_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14665_ net1378 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__inv_2
X_11877_ net2070 net262 net484 vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16404_ clknet_leaf_77_wb_clk_i net1968 _00387_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09076__A0 _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13616_ net187 _04055_ _04056_ net728 vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17384_ clknet_leaf_30_wb_clk_i _03071_ _01367_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10828_ _07060_ _07100_ net329 _07082_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14596_ net1333 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__inv_2
XANTENNA__09615__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16335_ clknet_leaf_67_wb_clk_i _02089_ _00318_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_13547_ net185 _03997_ _03998_ net725 vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__a211o_1
X_10759_ net528 _06935_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__nor2_2
XFILLER_0_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09629__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16266_ clknet_leaf_107_wb_clk_i net1720 _00254_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
XANTENNA__17033__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13478_ _03934_ _03936_ _03938_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18005_ net1505 vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_hd__buf_2
XFILLER_0_129_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13175__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15217_ net1292 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12429_ net3155 net247 net416 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16197_ clknet_leaf_115_wb_clk_i _01957_ _00185_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10918__D1 _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13580__C1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15148_ net1197 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10933__A1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07970_ net1062 vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__inv_2
X_15079_ net1300 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18070__1570 vssd1 vssd1 vccd1 vccd1 _18070__1570/HI net1570 sky130_fd_sc_hd__conb_1
XFILLER_0_120_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08354__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[23\] net966
+ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_69_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_109_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09571_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[25\] net971
+ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_65_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08522_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[18\] net882
+ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__and3_1
XANTENNA__11833__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08708__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08453_ net1106 net1112 net1115 net1109 vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_4_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08384_ net729 net720 vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14060__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08814__B1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12664__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout417_A _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1061_A team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14445__A net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1159_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10621__B1 _06960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08443__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09005_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[9\] net908 vssd1
+ vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13166__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11177__A1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17526__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1326_A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08042__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout786_A _04659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__A1 _04969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08593__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout510 _05996_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout521 net522 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09907_ _06234_ _06235_ _06245_ _06246_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__or4_1
Xfanout532 _05222_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_2
XANTENNA__16550__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17676__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout543 net544 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_4
Xfanout554 net555 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09705__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout953_A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 _04620_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__buf_2
XFILLER_0_77_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout576 _07792_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__dlymetal6s2s_1
X_09838_ _06167_ _06170_ _06172_ _06177_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__or4_1
Xfanout587 net590 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_4
Xfanout598 net599 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__buf_4
XANTENNA__10152__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12839__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[15\] net803 net754 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ net3131 net207 net491 vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[16\] _07541_ net1028 vssd1 vssd1
+ vccd1 vccd1 _03615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11731_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[5\] net718 vssd1 vssd1 vccd1
+ vccd1 _07922_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14450_ net1374 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11662_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[19\] _07135_ net716 vssd1 vssd1
+ vccd1 vccd1 _07867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14051__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13401_ _03860_ _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__nand2b_1
X_10613_ _06951_ _06952_ vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_94_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12574__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14381_ net1316 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11593_ _07809_ vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__inv_2
X_16120_ clknet_leaf_101_wb_clk_i _01895_ _00108_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13332_ net564 _07702_ _03808_ net585 vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10544_ _05805_ _05807_ _05835_ net560 vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__a31o_1
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire955 net956 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_126_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16051_ clknet_leaf_87_wb_clk_i _01844_ _00039_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13263_ net1062 _03754_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1
+ vccd1 _03755_ sky130_fd_sc_hd__o21ai_1
X_10475_ net504 _06780_ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15002_ net1190 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12214_ net3272 net303 net444 vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13194_ net15 net837 net630 net3213 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__a22o_1
XANTENNA__08033__B2 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10915__A1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11918__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15186__A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12145_ net2788 net228 net452 vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_7_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_88_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10391__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13314__C1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12076_ net2190 net261 net460 vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__mux2_1
X_16953_ clknet_leaf_51_wb_clk_i _02640_ _00936_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15904_ net1336 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__inv_2
X_11027_ _05491_ _06158_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__xor2_1
XANTENNA__10679__B1 _07018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16884_ clknet_leaf_12_wb_clk_i _02571_ _00867_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10143__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15835_ net1373 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__inv_2
XANTENNA__13617__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11576__A_N team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13093__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15766_ net1346 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12978_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[108\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[116\]
+ net858 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__mux2_1
XANTENNA__08528__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09836__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17505_ clknet_leaf_48_wb_clk_i _03192_ _01488_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14717_ net1309 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11929_ net2844 net219 net477 vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__mux2_1
XANTENNA__12840__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15697_ net1341 vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10496__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17436_ clknet_leaf_37_wb_clk_i _03123_ _01419_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14648_ net1180 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_70_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_111_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14042__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_17 _06737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 _07873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12484__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ clknet_leaf_128_wb_clk_i _03054_ _01350_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14579_ net1408 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__inv_2
XANTENNA__16423__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17549__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16318_ clknet_leaf_68_wb_clk_i _02072_ _00301_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08272__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17298_ clknet_leaf_129_wb_clk_i _02985_ _01281_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16249_ clknet_leaf_107_wb_clk_i net1793 _00237_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11159__A1 _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
XANTENNA__11159__B2 _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_3_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13553__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_88_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17699__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_120_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XANTENNA__11828__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
Xoutput179 net636 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09094__A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11331__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10765__S0 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09623_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] net625 _05961_ _05962_
+ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__a22o_2
XFILLER_0_78_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12659__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13608__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09554_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[28\] net816 net738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17079__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09827__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08505_ net730 _04752_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1
+ vccd1 vccd1 _04845_ sky130_fd_sc_hd__o21a_1
XANTENNA__12831__A1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09485_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[30\] net666 net657 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout534_A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1276_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08436_ net1013 net914 vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__and2_2
XFILLER_0_93_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14033__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_77_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12394__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08367_ _04706_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout701_A _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08298_ net1151 net1153 net1147 net1150 vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__and4bb_1
XANTENNA__09460__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16916__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13139__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10260_ _06133_ _06162_ _06165_ _06599_ _06132_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__o221a_1
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10191_ _06528_ _06529_ _06526_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10642__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_115_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1305 net1306 vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__buf_4
XFILLER_0_44_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1316 net1317 vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__buf_4
XFILLER_0_100_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1327 net1329 vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__buf_4
Xfanout1338 net1339 vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__buf_4
Xfanout340 _06590_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_4
Xfanout1349 net1351 vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__buf_4
Xfanout351 net352 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__buf_2
Xfanout362 _03653_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_2
X_13950_ _04223_ _04227_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__nand2_2
Xfanout373 _06465_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_2
Xfanout384 _03570_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_4
Xfanout395 _03567_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_8
X_12901_ net361 _03675_ net1029 vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13881_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[3\] _04187_ vssd1 vssd1 vccd1
+ vccd1 _04188_ sky130_fd_sc_hd__and2_1
XANTENNA__12569__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15620_ net1193 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__inv_2
XANTENNA__13254__A team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_57_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12832_ net1830 net640 net607 _03650_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__a22o_1
XANTENNA__08348__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15551_ net1256 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12763_ net2025 net642 net609 _03603_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14502_ net1335 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__inv_2
X_11714_ net3012 net284 net502 vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15482_ net1193 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__inv_2
XANTENNA__14024__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12694_ net3253 net212 net385 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__mux2_1
X_17221_ clknet_leaf_40_wb_clk_i _02908_ _01204_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14433_ net1381 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__inv_2
X_11645_ _07817_ _07853_ vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__and2b_1
X_17152_ clknet_leaf_33_wb_clk_i _02839_ _01135_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09179__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_14364_ net1352 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11576_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\]
+ vssd1 vssd1 vccd1 vccd1 _07793_ sky130_fd_sc_hd__and2b_2
Xinput37 gpio_in[19] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
XFILLER_0_135_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput48 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
X_16103_ clknet_leaf_92_wb_clk_i _01878_ _00091_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13315_ _04475_ _07706_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__nand2_1
XANTENNA__08514__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput59 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
X_17083_ clknet_leaf_17_wb_clk_i _02770_ _01066_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10527_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[31\] _04766_ net673
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[31\] _06866_ vssd1 vssd1 vccd1
+ vccd1 _06867_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14295_ net1355 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16034_ clknet_leaf_103_wb_clk_i net1663 _00028_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10458_ _06795_ _06796_ _06797_ vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__or3_1
X_13246_ net2186 net355 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1
+ vccd1 vccd1 _01904_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12889__A1 _05704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11648__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10552__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13429__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10389_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[16\] net816 _06727_
+ _06728_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__a211o_1
X_13177_ net1 _03732_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12128_ net2756 net218 net451 vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__mux2_1
X_17985_ net1485 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
XANTENNA__09345__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13302__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16936_ clknet_leaf_30_wb_clk_i _02623_ _00919_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15644__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12059_ net2732 net189 net459 vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__mux2_1
XANTENNA__10116__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11313__A1 _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17221__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12479__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16867_ clknet_leaf_22_wb_clk_i _02554_ _00850_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15818_ net1310 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__inv_2
X_16798_ clknet_leaf_46_wb_clk_i _02485_ _00781_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09080__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15749_ net1401 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__inv_2
XANTENNA__17371__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09270_ _05604_ _05605_ _05607_ _05609_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14015__B1 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08221_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[60\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[52\]
+ net1041 vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__mux2_1
X_17419_ clknet_leaf_1_wb_clk_i _03106_ _01402_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10727__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09089__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08152_ net829 net564 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09442__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08424__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08083_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[2\] net569 _04525_ _04556_
+ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__a22o_1
XANTENNA__15819__A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13541__A2 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_124_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_122_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1024_A _04490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__B net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[8\] net925 vssd1
+ vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout484_A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10107__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12389__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1393_A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16469__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_A _04682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08720__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09606_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[24\] net946
+ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11068__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09537_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[28\] net973 vssd1
+ vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__and3_1
XANTENNA__12804__A1 _07290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout916_A net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14006__B1 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09468_ net560 _05805_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__o21a_1
XANTENNA__09681__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08419_ net1107 net1114 net1113 net1110 vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__and4bb_4
X_09399_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[27\] net692 net666 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__a22o_1
XANTENNA__13013__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11430_ team_01_WB.instance_to_wrap.cpu.f0.i\[11\] _07676_ net610 team_01_WB.instance_to_wrap.cpu.f0.i\[12\]
+ vssd1 vssd1 vccd1 vccd1 _07740_ sky130_fd_sc_hd__a31o_1
XANTENNA__09433__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14055__D _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11361_ team_01_WB.instance_to_wrap.cpu.f0.i\[16\] team_01_WB.instance_to_wrap.cpu.f0.i\[15\]
+ _07689_ vssd1 vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__and3_1
XANTENNA__11240__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12852__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15729__A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13517__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10312_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[18\] net782 net740 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__a22o_1
X_13100_ net52 net51 net54 net53 vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__or4_1
XFILLER_0_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14080_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[100\] _04244_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[116\]
+ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__a22o_1
X_11292_ _07628_ net1155 _07631_ vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__mux2_1
XANTENNA__08631__A team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08539__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10243_ _06576_ _06577_ _06578_ _06582_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__or4_1
X_13031_ net2461 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[63\] net861 vssd1 vssd1
+ vccd1 vccd1 _02094_ sky130_fd_sc_hd__mux2_1
XANTENNA__11543__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12740__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17244__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[10\] net812 net757 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__a22o_1
Xfanout1102 net1104 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input45_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1113 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[21\] vssd1 vssd1 vccd1 vccd1
+ net1113 sky130_fd_sc_hd__clkbuf_2
Xfanout1124 net1126 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__buf_2
Xfanout1135 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1 vccd1 vccd1
+ net1135 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15464__A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17770_ clknet_leaf_76_wb_clk_i _03446_ _01710_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[40\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1146 net1147 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__clkbuf_2
X_14982_ net1299 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__inv_2
Xfanout1157 team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1 net1157
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13296__A1 _07650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10104__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1179 net1182 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__buf_2
Xfanout192 _07823_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_2
X_16721_ clknet_leaf_14_wb_clk_i _02408_ _00704_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13933_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__nand2_8
XANTENNA__12299__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17394__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16652_ clknet_leaf_133_wb_clk_i _02339_ _00635_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13864_ net1164 net1058 net3284 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[25\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_9_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10401__A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15603_ net1279 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08509__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12815_ net1033 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[5\] vssd1 vssd1 vccd1
+ vccd1 _03639_ sky130_fd_sc_hd__or2_1
X_16583_ clknet_leaf_123_wb_clk_i _02270_ _00566_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13795_ _04165_ _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11931__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15534_ net1283 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ net3203 net639 net606 _03591_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15465_ net1230 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__inv_2
X_12677_ net2464 net284 net388 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17204_ clknet_leaf_13_wb_clk_i _02891_ _01187_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14416_ net1348 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__inv_2
X_11628_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _07818_ vssd1 vssd1
+ vccd1 vccd1 _07840_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15396_ net1191 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__inv_2
XANTENNA__09424__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17135_ clknet_leaf_141_wb_clk_i _02822_ _01118_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13771__A2 _04152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09975__B2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15639__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14347_ net1370 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__inv_2
X_11559_ _07787_ _07788_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire582 _06517_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10585__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[14\] vssd1 vssd1 vccd1 vccd1
+ net2234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold629 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[90\] vssd1 vssd1 vccd1 vccd1
+ net2245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09637__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17066_ clknet_leaf_11_wb_clk_i _02753_ _01049_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14278_ net1367 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09727__A1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16017_ net1386 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__inv_2
X_13229_ net2877 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1
+ vccd1 vccd1 _01921_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11534__B2 net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1307 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2923 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08950__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_6__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__16611__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08770_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] net702 _05104_ _05109_
+ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__o22a_4
Xhold1318 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2934 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13287__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17968_ net1468 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1329 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16919_ clknet_leaf_138_wb_clk_i _02606_ _00902_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_17899_ net1419 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08702__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12002__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11841__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09322_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[24\] net681 net670 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08716__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09253_ net600 _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17117__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout232_A net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08204_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[77\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[69\]
+ net1039 vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09184_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[16\] net879
+ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08135_ _04489_ team_01_WB.instance_to_wrap.cpu.f0.num\[0\] team_01_WB.instance_to_wrap.cpu.f0.num\[19\]
+ _04475_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_71_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12672__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1141_A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10576__A2 _06882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11773__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1239_A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ _04512_ _04529_ _04539_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__a21oi_1
XANTENNA__17267__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout699_A _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13514__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1406_A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11525__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout866_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08968_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[8\] net896 vssd1
+ vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_51_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09282__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08899_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[2\] net887 vssd1
+ vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10930_ _06469_ _06472_ _06568_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_92_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10861_ net525 _07123_ _07149_ _06957_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_21_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12847__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12600_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[20\] net272 net397 vssd1
+ vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13580_ net200 net196 _07879_ net646 vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10792_ net515 _06897_ _07120_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__o21a_1
XANTENNA__13450__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12531_ net3023 net206 net403 vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08345__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14066__C _04348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15250_ net1232 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__inv_2
XANTENNA__09406__B1 _04797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12462_ net3055 net247 net413 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14201_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\] vssd1 vssd1 vccd1
+ vccd1 _02286_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11413_ _07693_ _07729_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15181_ net1215 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__inv_2
XANTENNA__12582__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12393_ net2492 net222 net419 vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__mux2_1
XANTENNA__11202__D _07541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12961__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14132_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[71\] _04247_ _04249_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11344_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\] team_01_WB.instance_to_wrap.cpu.f0.i\[1\]
+ _07671_ vssd1 vssd1 vccd1 vccd1 _07673_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16634__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14063_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[99\] _04254_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[123\]
+ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__a22o_1
X_11275_ _07038_ _07100_ net329 _07029_ vssd1 vssd1 vccd1 vccd1 _07615_ sky130_fd_sc_hd__a22o_1
XANTENNA__11516__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10319__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13014_ net2303 net1633 net868 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__mux2_1
X_10226_ _06562_ _06565_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__nand2_1
XANTENNA__11926__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17822_ clknet_leaf_64_wb_clk_i _03498_ _01762_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[92\]
+ sky130_fd_sc_hd__dfstp_1
X_10157_ net561 _04970_ net343 vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__or3_1
XANTENNA__13269__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_101_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4 _01985_ vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09192__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16784__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14965_ net1225 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__inv_2
X_17753_ clknet_leaf_79_wb_clk_i net3016 _01693_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10088_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[7\] net761 _06417_ _06420_
+ net768 vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_106_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13916_ _04142_ _04207_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__and2_1
X_16704_ clknet_leaf_29_wb_clk_i _02391_ _00687_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15922__A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10131__A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17684_ clknet_leaf_94_wb_clk_i _03368_ _01625_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_102_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14896_ net1223 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
X_17949__1449 vssd1 vssd1 vccd1 vccd1 _17949__1449/HI net1449 sky130_fd_sc_hd__conb_1
X_16635_ clknet_leaf_50_wb_clk_i _02322_ _00618_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13847_ net1166 net1060 net2424 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[8\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_58_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11661__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13442__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16566_ clknet_leaf_109_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_dhit _00549_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.dhit sky130_fd_sc_hd__dfrtp_2
X_13778_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[2\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ net604 vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09645__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15517_ net1252 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_119_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12729_ _03575_ _03578_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13992__A2 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16497_ clknet_leaf_106_wb_clk_i _02251_ _00480_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16164__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15448_ net1195 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15369__A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12492__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15379_ net1278 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12952__A0 team_01_WB.instance_to_wrap.cpu.f0.write_data\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17118_ clknet_leaf_44_wb_clk_i _02805_ _01101_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold404 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold415 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[23\] vssd1 vssd1 vccd1 vccd1 net2031
+ sky130_fd_sc_hd__dlygate4sd3_1
X_18098_ net637 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_1
Xhold426 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14154__C1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold448 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] net627 _06278_ _06279_
+ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__a22o_2
X_17049_ clknet_leaf_51_wb_clk_i _02736_ _01032_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout906 net907 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__clkbuf_4
X_09871_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[12\] net745 net737 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__a22o_1
Xfanout928 net929 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout939 _04756_ vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11836__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[1\] net937 vssd1
+ vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__and3_1
XANTENNA__10740__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10191__B1 _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2731 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2753 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net1088 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[4\] net901 vssd1
+ vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__and3_1
Xhold1148 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2764 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09533__C net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1159 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2775 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10041__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08684_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[7\] net885 vssd1
+ vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11691__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12667__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1091_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_A _07958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1189_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16507__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09305_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[22\] net679 _05630_
+ _05636_ _05637_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_130_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11443__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13983__A2 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10797__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1356_A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09236_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[21\] net668 _05574_ _05575_
+ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_131_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09939__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13196__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13735__A2 _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09167_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[16\] net881
+ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09403__A3 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12943__B1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11746__B2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11600__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09277__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08118_ net1063 _04495_ team_01_WB.instance_to_wrap.cpu.f0.num\[18\] _04476_ vssd1
+ vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__a22o_1
XANTENNA__08611__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[13\] net933 vssd1
+ vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout983_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09708__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08049_ _04521_ team_01_WB.instance_to_wrap.cpu.K0.code\[3\] team_01_WB.instance_to_wrap.cpu.K0.code\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_129_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold960 _03517_ vssd1 vssd1 vccd1 vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14911__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold971 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[33\] vssd1 vssd1 vccd1 vccd1
+ net2587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11060_ net373 _07380_ _05301_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__nor3b_1
Xhold982 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 _02113_ vssd1 vssd1 vccd1 vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10011_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[1\] net752 net771 vssd1
+ vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__a21o_1
XANTENNA__08914__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10182__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09443__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13120__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11047__A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1660 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14750_ net1309 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__inv_2
Xhold1671 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 net3287
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11962_ net2545 _07831_ net473 vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__mux2_1
XANTENNA__09875__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13701_ _04106_ _04119_ _04121_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[9\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_58_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10913_ _06596_ _07252_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12577__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14681_ net1343 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__inv_2
X_11893_ net2720 net190 net480 vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16420_ clknet_leaf_104_wb_clk_i _02174_ _00403_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13262__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13632_ net200 net196 _07911_ net646 vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__o211a_1
X_10844_ net339 _07016_ net330 _07183_ _07179_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__a221o_1
XANTENNA__16187__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13423__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13423__B2 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16351_ clknet_leaf_67_wb_clk_i _02105_ _00334_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13563_ net198 net194 _07869_ net643 vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10775_ _06675_ _07114_ _06641_ vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11985__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15302_ net1324 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12514_ net2251 net279 net407 vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16282_ clknet_leaf_63_wb_clk_i _02036_ _00265_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_114_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08850__A1 _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13494_ _03952_ _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_97_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18021_ net1521 vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_114_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13187__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15233_ net1248 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__inv_2
X_12445_ net2054 net252 net417 vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12934__B1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15164_ net1175 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__inv_2
X_12376_ net2439 net256 net425 vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14115_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[62\] _04260_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__a22o_1
XANTENNA__08522__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11327_ _07661_ net2047 _07655_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15095_ net1199 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09915__A _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output76_A net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[35\] _04221_ _04230_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[35\]
+ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__a22o_1
XANTENNA__14151__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11258_ _06966_ _07278_ _06964_ vssd1 vssd1 vccd1 vccd1 _07598_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08366__B1 _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11656__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10209_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[8\] net819 net812 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11189_ _06921_ _07527_ _07528_ _07185_ vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_66_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17805_ clknet_leaf_72_wb_clk_i net2868 _01745_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15997_ net1407 vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10499__C _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17736_ clknet_leaf_84_wb_clk_i net1961 _01676_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14948_ net1239 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__inv_2
XANTENNA__09866__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13662__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09330__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10476__A1 _05931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12487__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17667_ clknet_leaf_117_wb_clk_i _03352_ _01608_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14879_ net1256 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16618_ clknet_leaf_3_wb_clk_i _02305_ _00601_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17598_ clknet_leaf_69_wb_clk_i _03285_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09618__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16549_ clknet_leaf_111_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[15\]
+ _00532_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11404__B net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11976__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09021_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[9\] net924 vssd1
+ vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13178__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold201 team_01_WB.instance_to_wrap.cpu.f0.write_data\[23\] vssd1 vssd1 vccd1 vccd1
+ net1817 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold212 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 net113 vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold234 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 _01984_ vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[15\] vssd1 vssd1 vccd1 vccd1
+ net1894 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[4\] net965 vssd1
+ vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__and3_1
Xhold289 _02153_ vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout703 _04758_ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__buf_4
XANTENNA__14142__A2 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08357__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13853__A_N net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 net726 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout397_A _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout736 _04687_ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__buf_4
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09854_ _06192_ _06193_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__nand2b_1
Xfanout747 _04682_ vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__clkbuf_4
Xfanout758 _04675_ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_8
Xfanout769 _04672_ vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1104_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[0\] net892 vssd1
+ vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__and3_1
XANTENNA__11468__A1_N net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09785_ _06109_ _06110_ _06123_ _06124_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__or4_1
XFILLER_0_119_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15562__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08736_ net603 _05074_ _05075_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__a21o_2
XFILLER_0_59_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13653__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10202__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17455__CLK clknet_leaf_143_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09321__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout731_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12397__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[7\] net910 vssd1
+ vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18019__1519 vssd1 vssd1 vccd1 vccd1 _18019__1519/HI net1519 sky130_fd_sc_hd__conb_1
XFILLER_0_95_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09609__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[15\] net687 net666 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11314__B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10560_ _04741_ _04743_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__nand2_2
XFILLER_0_130_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13169__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[17\] net683 _05547_
+ _05548_ _05552_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_49_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10491_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[31\] net976
+ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12916__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ net2848 net214 net441 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11825__A_N team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08596__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12860__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15737__A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12161_ net2947 net217 net447 vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__mux2_1
X_17948__1448 vssd1 vssd1 vccd1 vccd1 _17948__1448/HI net1448 sky130_fd_sc_hd__conb_1
XANTENNA__14641__A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10942__A2 _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11112_ net550 net373 _06946_ vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_102_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14133__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12092_ net3158 net189 net455 vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold790 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13257__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ _05076_ _06250_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__nand2_1
X_15920_ net1330 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__inv_2
XANTENNA__10155__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15851_ net1364 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09173__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14802_ net1228 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15782_ net1307 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__inv_2
X_12994_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[92\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[100\]
+ net858 vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__mux2_1
XANTENNA__09848__B1 _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13644__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09470__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1490 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3106 sky130_fd_sc_hd__dlygate4sd3_1
X_14733_ net1319 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__inv_2
XANTENNA__09312__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17521_ clknet_leaf_14_wb_clk_i _03208_ _01504_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11945_ net1903 net290 net477 vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17452_ clknet_leaf_134_wb_clk_i _03139_ _01435_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16822__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11505__A team_01_WB.instance_to_wrap.cpu.DM0.data_i\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14664_ net1382 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__inv_2
XANTENNA__12100__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11876_ net2335 net233 net485 vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ clknet_leaf_86_wb_clk_i net1941 _00386_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08517__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13615_ net199 net195 _07806_ _07899_ net645 vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__o2111a_1
XANTENNA__09076__A1 _05415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17383_ clknet_leaf_16_wb_clk_i _03070_ _01366_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10827_ net370 _07165_ _07166_ net507 _05619_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__o32a_1
X_14595_ net1392 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16334_ clknet_leaf_68_wb_clk_i net2787 _00317_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13546_ net197 net193 _07857_ net643 vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__o211a_1
X_10758_ _04844_ net332 _07094_ net370 _07097_ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16265_ clknet_leaf_106_wb_clk_i net1917 _00253_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13477_ _04500_ _04842_ _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10689_ _07027_ _07028_ net517 vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_33_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18004_ net1504 vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_hd__buf_2
X_15216_ net1271 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12428_ net3267 net214 net416 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__mux2_1
XANTENNA__09379__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16196_ clknet_leaf_115_wb_clk_i _01956_ _00184_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10918__C1 _05374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14109__C1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15147_ net1297 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16202__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12359_ net2874 net223 net423 vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17328__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14124__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15078_ net1292 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__inv_2
X_14029_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] _04249_ _04259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[18\]
+ _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__a221o_1
XANTENNA__09551__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09083__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09570_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[25\] net950 vssd1
+ vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__and3_1
XANTENNA__09839__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13635__A1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08521_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[18\] net931
+ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__and3_1
X_17719_ clknet_leaf_109_wb_clk_i _00014_ _01660_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_77_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11415__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12010__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[23\] net938
+ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_19_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08383_ net1156 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\]
+ _04711_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__or4_4
XFILLER_0_110_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10973__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout312_A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08443__B net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1054_A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09004_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[9\] net916 vssd1
+ vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11150__A _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15557__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12680__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1221_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14461__A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08042__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_105_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_44_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14115__A2 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout681_A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout500 _07795_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout779_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 _05963_ vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13323__B1 _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout522 _05260_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_2
X_09906_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[5\] net817 net753 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout533 net536 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10137__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__buf_2
Xfanout555 _05114_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_2
Xfanout566 _04620_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_1
X_09837_ _06173_ _06174_ _06175_ _06176_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__or4_1
Xfanout577 _07753_ vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_2
Xfanout588 net590 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout599 _04755_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout946_A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16845__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13626__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[15\] net751 net742 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09290__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08719_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[5\] net890 vssd1
+ vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09699_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[21\] net948 vssd1
+ vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_29_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08502__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11730_ net2641 net300 net502 vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16995__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08337__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11661_ net1990 net273 net500 vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__mux2_1
XANTENNA__12855__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] net595 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__a21o_1
X_10612_ net550 _06339_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14380_ net1319 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11592_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] _07808_ vssd1 vssd1
+ vccd1 vccd1 _07809_ sky130_fd_sc_hd__and2_2
XANTENNA__08634__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10883__B _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_144_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_52_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13331_ _04479_ _07686_ _03743_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__a21oi_1
XANTENNA__16225__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10543_ net503 _06882_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__xor2_2
XFILLER_0_134_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire956 _04656_ vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11060__A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16050_ clknet_leaf_87_wb_clk_i _01843_ _00038_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13262_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] _03753_ vssd1 vssd1 vccd1 vccd1
+ _03754_ sky130_fd_sc_hd__or2_1
X_10474_ _06811_ _06813_ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__and2_1
XANTENNA__09168__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15001_ net1258 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__inv_2
X_12213_ net2687 net284 net446 vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12590__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13193_ net16 net835 net628 net3039 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__o22a_1
XANTENNA__08033__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10915__A2 _06738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14106__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12144_ net2598 net287 net452 vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__mux2_1
XANTENNA__09781__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16952_ clknet_leaf_27_wb_clk_i _02639_ _00935_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12075_ net3225 net231 net461 vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__mux2_1
X_15903_ net1409 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__inv_2
X_11026_ _04947_ net375 vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__xor2_1
XANTENNA__10679__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16883_ clknet_leaf_135_wb_clk_i _02570_ _00866_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11934__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15834_ net1372 vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13617__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12977_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[109\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[117\]
+ net857 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__mux2_1
XANTENNA__09631__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15765_ net1346 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17504_ clknet_leaf_29_wb_clk_i _03191_ _01487_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15930__A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14716_ net1309 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__inv_2
X_11928_ net2799 net220 net477 vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__mux2_1
X_15696_ net1224 vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17000__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17435_ clknet_leaf_20_wb_clk_i _03122_ _01418_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14647_ net1188 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11859_ net575 _07793_ _07946_ vssd1 vssd1 vccd1 vccd1 _07948_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_18 _07827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14578_ net1388 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__inv_2
X_17366_ clknet_leaf_1_wb_clk_i _03053_ _01349_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_29 _07873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16317_ clknet_leaf_75_wb_clk_i _02071_ _00300_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_13529_ net186 _03982_ _03983_ net726 vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__a211o_1
X_17297_ clknet_leaf_14_wb_clk_i _02984_ _01280_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16248_ clknet_leaf_95_wb_clk_i _02008_ _00236_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_2_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
X_16179_ clknet_leaf_107_wb_clk_i _01939_ _00167_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10367__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XANTENNA__10906__A2 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09772__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
X_18018__1518 vssd1 vssd1 vccd1 vccd1 _18018__1518/HI net1518 sky130_fd_sc_hd__conb_1
XANTENNA__08710__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12005__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10119__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10314__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11844__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11331__A2 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] net764 net622 vssd1
+ vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__o21a_1
XANTENNA__10765__S1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13608__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08719__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11619__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _05876_ _05890_ _05891_ _05892_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__or4_1
XANTENNA__09541__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout262_A _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08438__B net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11145__A _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08504_ net598 _04837_ _04843_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__o21a_2
X_09484_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[30\] net647 _05812_
+ _05813_ _05815_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__a2111o_1
X_17947__1447 vssd1 vssd1 vccd1 vccd1 _17947__1447/HI net1447 sky130_fd_sc_hd__conb_1
XFILLER_0_77_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08435_ net1107 net1110 net1112 net1114 vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__nor4b_1
XANTENNA__12675__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1171_A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13360__A team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1269_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08366_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] net625 _04704_ _04705_
+ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__a22o_4
XFILLER_0_46_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08454__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08297_ net988 net975 vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16398__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17643__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout896_A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10923__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10358__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09285__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ _06526_ _06528_ _06529_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1306 net1314 vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__buf_4
Xfanout1317 net1322 vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__buf_4
Xfanout1328 net1329 vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__clkbuf_4
Xfanout330 _07070_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_4
Xfanout1339 net1340 vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__buf_4
Xfanout341 _06495_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_4
Xfanout352 _03742_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout363 net364 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_2
Xfanout374 _06188_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_2
Xfanout385 _03570_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_6
Xfanout396 _03567_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_4
X_12900_ _05654_ net577 vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__nor2_1
X_13880_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[2\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[1\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _04187_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_134_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12831_ net1034 _07438_ net366 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\]
+ net1057 vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__a32o_1
XFILLER_0_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08348__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15550_ net1248 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12762_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] net1055 net363 _03602_
+ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14501_ net1398 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11713_ net612 _07802_ _07907_ _07906_ vssd1 vssd1 vccd1 vccd1 _07908_ sky130_fd_sc_hd__a31o_4
XFILLER_0_16_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15481_ net1260 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12585__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12693_ net2956 net247 net385 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14432_ net1381 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__inv_2
X_17220_ clknet_leaf_53_wb_clk_i _02907_ _01203_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11644_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\]
+ _07814_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1 vccd1 vccd1
+ _07853_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17151_ clknet_leaf_26_wb_clk_i _02838_ _01134_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14363_ net1352 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10597__A0 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
X_11575_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] _07784_ _07789_ vssd1 vssd1
+ vccd1 vccd1 _07792_ sky130_fd_sc_hd__and3_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16102_ clknet_leaf_91_wb_clk_i _01877_ _00090_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput38 wb_rst_i vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
X_13314_ _07686_ _07708_ _03794_ net586 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__o211a_1
X_17082_ clknet_leaf_45_wb_clk_i _02769_ _01065_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10526_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[31\] net677 net666 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__a22o_1
Xinput49 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14294_ net1355 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16033_ clknet_leaf_106_wb_clk_i _01827_ _00027_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13535__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11929__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15197__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13245_ net2750 net356 net352 team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1
+ vccd1 vccd1 _01905_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10457_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[26\] net787 net752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09195__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09754__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ net108 net850 net842 net2015 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a22o_1
XANTENNA__13429__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10388_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[16\] net810 net774 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08530__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12127_ net2364 net221 net454 vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_5__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_17984_ net1484 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XANTENNA__10134__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12058_ _07790_ net576 _07951_ vssd1 vssd1 vccd1 vccd1 _07955_ sky130_fd_sc_hd__and3_4
XFILLER_0_40_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16935_ clknet_leaf_15_wb_clk_i _02622_ _00918_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13445__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ _05707_ net512 vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__xnor2_1
X_16866_ clknet_leaf_34_wb_clk_i _02553_ _00849_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_15817_ net1311 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__inv_2
X_16797_ clknet_leaf_20_wb_clk_i _02484_ _00780_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17516__CLK clknet_leaf_132_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15748_ net1240 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12813__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12495__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14015__B2 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08493__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15679_ net1260 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__inv_2
X_08220_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[61\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[53\]
+ net1039 vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17418_ clknet_leaf_2_wb_clk_i _03105_ _01401_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08705__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08151_ net564 vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__inv_2
XANTENNA__11234__D1 _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17349_ clknet_leaf_38_wb_clk_i _03036_ _01332_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09442__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10309__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10052__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08082_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\] _04555_ _04524_ vssd1 vssd1 vccd1
+ vccd1 _04556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12329__A1 _07838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11839__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16690__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09745__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11552__A2 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08984_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[8\] net671 _05321_ _05322_
+ _05323_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1017_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17046__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12501__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08449__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10512__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09605_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[24\] net964 vssd1
+ vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17196__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1386_A net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[28\] net790 net741 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11068__B2 _05374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09467_ _05760_ _05781_ net378 vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout811_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout909_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08418_ net1004 net938 vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__nand2_4
XANTENNA__11603__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09398_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\] net699 net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[30\] net964 vssd1
+ vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10043__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11360_ net1065 _07676_ _07682_ vssd1 vssd1 vccd1 vccd1 _07689_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11749__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[18\] net811 net800 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11291_ _06886_ _06887_ _06960_ _04492_ vssd1 vssd1 vccd1 vccd1 _07631_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08631__B net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13030_ net1933 net1874 net868 vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__mux2_1
X_10242_ _06571_ _06579_ _06580_ _06581_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__or4_1
XANTENNA__14190__B1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09446__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12740__B2 _03587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15745__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ _06509_ _06510_ _06511_ _06512_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__or4_1
Xfanout1103 net1104 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1114 net1115 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_2
Xfanout1125 net1126 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__buf_1
Xfanout1136 net1137 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input38_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1 vccd1
+ net1147 sky130_fd_sc_hd__clkbuf_2
X_14981_ net1206 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__inv_2
Xfanout1158 net1160 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__buf_2
Xfanout1169 net1170 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__buf_2
X_16720_ clknet_leaf_127_wb_clk_i _02407_ _00703_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13932_ _04222_ _04223_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__nand2_2
Xfanout193 net194 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10503__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13863_ net1163 net1058 net2198 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[24\]
+ sky130_fd_sc_hd__and3b_1
X_16651_ clknet_leaf_4_wb_clk_i _02338_ _00634_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09181__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15602_ net1233 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
X_12814_ net1033 _07507_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13794_ _04160_ _04162_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__nor2_1
X_16582_ clknet_leaf_41_wb_clk_i _02269_ _00565_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16563__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15533_ net1215 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__inv_2
X_12745_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] net1054 net363 _03590_
+ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18017__1517 vssd1 vssd1 vccd1 vccd1 _18017__1517/HI net1517 sky130_fd_sc_hd__conb_1
XFILLER_0_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15464_ net1277 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__inv_2
XANTENNA__11096__A_N _07364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10282__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12676_ net2075 net251 net387 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17203_ clknet_leaf_135_wb_clk_i _02890_ _01186_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14415_ net1366 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__inv_2
XANTENNA__08525__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11627_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[26\] _07588_ net715 vssd1 vssd1
+ vccd1 vccd1 _07839_ sky130_fd_sc_hd__mux2_1
X_15395_ net1175 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_7_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14346_ net1375 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__inv_2
X_17134_ clknet_leaf_8_wb_clk_i _02821_ _01117_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11558_ team_01_WB.instance_to_wrap.cpu.K0.enable _07786_ net3277 vssd1 vssd1 vccd1
+ vccd1 _07788_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08822__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold608 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13508__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire583 _05040_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_4
X_10509_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[31\] net735 _06831_ _06836_
+ _06839_ vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__a2111o_1
X_17065_ clknet_leaf_10_wb_clk_i _02752_ _01048_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold619 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
X_14277_ net1368 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11489_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[18\] net579 vssd1 vssd1 vccd1
+ vccd1 _07772_ sky130_fd_sc_hd__nand2_1
XANTENNA__17069__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16016_ net1373 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__inv_2
X_13228_ net2114 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[22\] vssd1 vssd1
+ vccd1 vccd1 _01922_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17946__1446 vssd1 vssd1 vccd1 vccd1 _17946__1446/HI net1446 sky130_fd_sc_hd__conb_1
XANTENNA__11534__A2 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12731__A1 _06961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13159_ net1835 net843 net840 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[17\] vssd1
+ vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17967_ net1467 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
Xhold1308 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1319 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16918_ clknet_leaf_141_wb_clk_i _02605_ _00901_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17898_ net1418 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16906__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XANTENNA__09091__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16849_ clknet_leaf_18_wb_clk_i _02536_ _00832_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10030__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09321_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[24\] net657 net654 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[24\]
+ _05660_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12798__A1 _07531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09252_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[21\] net713 net594 vssd1 vssd1
+ vccd1 vccd1 _05592_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08203_ net2909 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[70\] net1042 vssd1 vssd1
+ vccd1 vccd1 _03484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09183_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[16\] net881 vssd1
+ vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10039__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13211__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10025__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08134_ _04600_ _04601_ _04602_ _04603_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_133_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09966__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08623__C1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08065_ _04538_ _04540_ _04541_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08451__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1134_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09718__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16436__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1301_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10205__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09563__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[8\] net667 _05304_ _05305_
+ _05306_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_127_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout761_A _04674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08898_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[2\] net890 vssd1
+ vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_123_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16586__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17831__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10860_ _07198_ _07199_ net519 vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12789__A1 _07553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13986__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09519_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[29\] net799 net792 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10791_ _07100_ _07123_ _07124_ net329 _07130_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12530_ net2812 net276 net405 vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_61_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11052__B _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12461_ net3163 net214 net413 vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__mux2_1
XANTENNA__12863__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13202__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14200_ _04154_ _04464_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_10_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10016__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11213__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11412_ team_01_WB.instance_to_wrap.cpu.f0.i\[19\] _07692_ net325 vssd1 vssd1 vccd1
+ vccd1 _07729_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15180_ net1180 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__inv_2
X_12392_ net2984 net223 net419 vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17211__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14131_ _04342_ _04396_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11343_ team_01_WB.instance_to_wrap.cpu.f0.i\[1\] _07671_ vssd1 vssd1 vccd1 vccd1
+ _07672_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14062_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[83\] _04245_ _04247_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[67\]
+ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__a221o_1
XANTENNA__09709__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11274_ net555 _07498_ vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__or2_1
XANTENNA__09176__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13013_ net3081 net2893 net867 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__mux2_1
XANTENNA__15475__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10225_ _05338_ _06564_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17821_ clknet_leaf_71_wb_clk_i net2352 _01761_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09473__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09590__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ net341 vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__inv_2
XANTENNA__13269__A2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5 team_01_WB.instance_to_wrap.a1.ADR_I\[20\] vssd1 vssd1 vccd1 vccd1 net1621
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17752_ clknet_leaf_86_wb_clk_i _03428_ _01692_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12103__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10412__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14964_ net1263 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__inv_2
X_10087_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[7\] net740 _06413_ _06414_
+ _06415_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_106_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08089__A _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16703_ clknet_leaf_26_wb_clk_i _02390_ _00686_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13915_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] _04185_ _04204_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17683_ clknet_leaf_81_wb_clk_i _03367_ _01624_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_14895_ net1214 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11942__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16634_ clknet_leaf_46_wb_clk_i _02321_ _00617_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13846_ net1167 net1060 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[7\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[7\] sky130_fd_sc_hd__and3b_1
XFILLER_0_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13977__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13442__B _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13777_ _04162_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__inv_2
X_16565_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[31\]
+ _00548_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10989_ _07005_ _07007_ vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15516_ net1172 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12728_ _04510_ _03578_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16496_ clknet_leaf_108_wb_clk_i _02250_ _00479_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12659_ net2961 net215 net389 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__mux2_1
X_15447_ net1195 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10007__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15378_ net1225 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08552__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12952__A1 _05300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17117_ clknet_leaf_40_wb_clk_i _02804_ _01100_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14329_ net1349 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__inv_2
Xhold405 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08620__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18097_ net637 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17704__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold427 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold438 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14154__B1 _04437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17048_ clknet_leaf_27_wb_clk_i _02735_ _01031_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold449 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[18\] vssd1 vssd1 vccd1 vccd1 net2065
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09086__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09870_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[12\] net805 net786 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__a22o_1
Xfanout907 net908 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__buf_4
XFILLER_0_1_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08821_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[1\] net927 vssd1
+ vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__and3_1
XANTENNA__17854__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1105 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\] vssd1 vssd1 vccd1 vccd1
+ net2721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1116 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2732 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[4\] net906 vssd1
+ vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__and3_1
Xhold1127 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2754 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12013__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10322__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1149 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2765 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08136__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09333__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11140__A0 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08683_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[7\] net915 vssd1
+ vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11852__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11691__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1084_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09304_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[22\] net651 _05623_ _05624_
+ _05633_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10246__A2 _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11443__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17234__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09235_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[21\] net665 net651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__a22o_1
XANTENNA__10797__A3 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12683__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout607_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1251_A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1349_A net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09939__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09166_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[16\] net896
+ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12943__A1 _05373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08117_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] team_01_WB.instance_to_wrap.cpu.f0.num\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11600__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09097_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[13\] net879
+ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17384__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_1__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14145__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08048_ net1774 net570 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[7\] vssd1 vssd1
+ vccd1 vccd1 _03543_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold950 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[18\] vssd1 vssd1 vccd1 vccd1
+ net2566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold961 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15295__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold983 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[98\] vssd1 vssd1 vccd1 vccd1
+ net2599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10010_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[1\] net801 net789 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_38_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09293__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18016__1516 vssd1 vssd1 vccd1 vccd1 _18016__1516/HI net1516 sky130_fd_sc_hd__conb_1
XFILLER_0_99_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09999_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] net627 _06337_ _06338_
+ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_34_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11636__A1_N net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3266 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09324__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11047__B _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1661 team_01_WB.instance_to_wrap.cpu.K0.count\[0\] vssd1 vssd1 vccd1 vccd1 net3277
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11961_ net2093 net225 net471 vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1672 team_01_WB.instance_to_wrap.cpu.c0.count\[13\] vssd1 vssd1 vccd1 vccd1 net3288
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12858__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11762__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10912_ _06469_ _06472_ _06568_ _06566_ vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__o31a_1
X_13700_ team_01_WB.instance_to_wrap.cpu.c0.count\[9\] _04105_ vssd1 vssd1 vccd1 vccd1
+ _04121_ sky130_fd_sc_hd__or2_1
X_14680_ net1365 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__inv_2
X_11892_ net575 _07942_ _07946_ vssd1 vssd1 vccd1 vccd1 _07949_ sky130_fd_sc_hd__and3_4
XFILLER_0_135_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_88_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13631_ _04051_ _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10843_ _07139_ _07182_ net524 vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17945__1445 vssd1 vssd1 vccd1 vccd1 _17945__1445/HI net1445 sky130_fd_sc_hd__conb_1
X_16350_ clknet_leaf_69_wb_clk_i _02104_ _00333_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10237__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13562_ _03921_ _03922_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10774_ _06712_ _06740_ _07112_ _06713_ _06677_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__a311o_1
XFILLER_0_66_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12513_ net3037 net303 net408 vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__mux2_1
X_15301_ net1210 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16281_ clknet_leaf_64_wb_clk_i _02035_ _00264_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12593__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13493_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] _03953_ vssd1 vssd1
+ vccd1 vccd1 _03954_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_97_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08850__A2 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16601__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18020_ net1520 vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_114_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12444_ net2846 net229 net417 vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__mux2_1
X_15232_ net1237 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08372__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08803__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12934__A1 _05415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15163_ net1180 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__inv_2
X_12375_ net2281 net260 net425 vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10945__A0 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14114_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[70\] _04233_ _04236_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[54\]
+ _04399_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__a221o_1
XANTENNA__14136__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11326_ _04548_ _07652_ _07660_ net1162 vssd1 vssd1 vccd1 vccd1 _07661_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15094_ net1202 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11937__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14045_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[91\] _04240_ _04243_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[27\]
+ _04333_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11257_ _07592_ _07593_ _07595_ _07596_ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__and4_1
XFILLER_0_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08366__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10208_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[8\] net824 _06535_ _06536_
+ _06544_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_108_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11188_ _06979_ _07240_ vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__nand2_1
XANTENNA__09634__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17107__CLK clknet_leaf_137_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17804_ clknet_leaf_66_wb_clk_i _03480_ _01744_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10139_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[11\] net798 net774 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15996_ net1387 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__inv_2
XANTENNA__08118__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13647__C1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17735_ clknet_leaf_85_wb_clk_i _03411_ _01675_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\]
+ sky130_fd_sc_hd__dfstp_1
X_14947_ net1187 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__inv_2
XANTENNA__14549__A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13662__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17666_ clknet_leaf_116_wb_clk_i _03351_ _01607_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14878_ net1274 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16617_ clknet_leaf_14_wb_clk_i _02304_ _00600_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13829_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[22\] net831 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[22\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_63_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17597_ clknet_leaf_69_wb_clk_i _03284_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10859__S0 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16548_ clknet_leaf_111_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[14\]
+ _00531_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16479_ clknet_leaf_92_wb_clk_i _02233_ _00462_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_116_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08841__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09020_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[9\] net908 vssd1
+ vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__and3_1
XANTENNA__13178__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12925__A1 _03692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08713__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold202 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12008__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09397__A3 _05707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold213 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[2\] vssd1 vssd1 vccd1 vccd1
+ net1829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _01980_ vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14127__B1 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold235 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 net1851
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold246 team_01_WB.instance_to_wrap.cpu.f0.write_data\[6\] vssd1 vssd1 vccd1 vccd1
+ net1862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11847__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold268 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09922_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[4\] net967 vssd1
+ vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout704 _04758_ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__buf_8
XFILLER_0_81_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout715 net716 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__clkbuf_4
Xfanout726 net729 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09554__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09853_ _06188_ _06191_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__nand2_1
Xfanout737 _04687_ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_124_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 _04682_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_6
XFILLER_0_42_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout292_A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout759 _04675_ vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_4
X_08804_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[0\] net675 _05141_ _05142_
+ _05143_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__a2111o_1
XANTENNA__15843__A net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[15\] net818 net801 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08735_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] net599 net596 vssd1 vssd1
+ vccd1 vccd1 _05075_ sky130_fd_sc_hd__and3_1
XANTENNA__12678__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1299_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08666_ _04971_ net584 net603 vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__mux2_2
XFILLER_0_90_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10467__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[15\] net939 net664 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[15\]
+ net707 vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_46_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10219__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_134_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09490__C1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09218_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[17\] net677 _05531_
+ _05539_ _05540_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_134_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09288__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10490_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[31\] net946
+ vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__and3_1
XANTENNA__16774__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12916__A1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09149_ _05480_ _05481_ _05487_ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_92_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08045__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10227__A _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14118__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12160_ net2581 net222 net448 vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ _06404_ _06405_ _07450_ vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__o21a_1
XANTENNA__10942__A3 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12091_ _07791_ net576 _07945_ vssd1 vssd1 vccd1 vccd1 _07956_ sky130_fd_sc_hd__and3_4
XFILLER_0_60_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold780 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[26\] vssd1 vssd1 vccd1 vccd1
+ net2396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09545__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11042_ _05076_ _06250_ vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10155__A1 _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15850_ net1363 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__inv_2
X_14801_ net1291 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__inv_2
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09848__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15781_ net1307 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__inv_2
X_12993_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[93\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[101\]
+ net857 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__mux2_1
XANTENNA__13644__A2 _07323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1480 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17520_ clknet_leaf_13_wb_clk_i _03207_ _01503_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1491 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3107 sky130_fd_sc_hd__dlygate4sd3_1
X_14732_ net1319 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__inv_2
XANTENNA__11655__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11944_ net2178 net257 net476 vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08367__A _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17451_ clknet_leaf_3_wb_clk_i _03138_ _01434_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11875_ net1910 net263 net484 vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__mux2_1
X_14663_ net1386 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__inv_2
XANTENNA_output107_A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ clknet_leaf_63_wb_clk_i _02156_ _00385_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[125\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_67_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13614_ _03887_ _04054_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__xnor2_1
X_10826_ net335 net337 _07164_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17382_ clknet_leaf_42_wb_clk_i _03069_ _01365_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14594_ net1401 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16333_ clknet_leaf_74_wb_clk_i _02087_ _00316_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13545_ _03928_ _03991_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__xnor2_1
X_10757_ _04844_ _05996_ net335 _07096_ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10091__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16264_ clknet_leaf_106_wb_clk_i net1920 _00252_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
X_13476_ _04500_ _04842_ _03927_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__o21ba_1
X_10688_ _06891_ _06937_ net533 vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09629__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18003_ net1503 vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_hd__buf_2
XFILLER_0_113_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12907__A1 _05615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15215_ net1213 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__inv_2
XANTENNA__08036__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12427_ net2374 net216 net415 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16195_ clknet_leaf_115_wb_clk_i _01955_ _00183_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13580__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09784__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15146_ net1276 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__inv_2
X_12358_ net3038 net190 net423 vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11667__S net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11309_ net727 _07438_ _07647_ vssd1 vssd1 vccd1 vccd1 _07648_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15077_ net1210 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12289_ net1952 net314 net438 vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14028_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[106\] _04252_ _04315_ _04317_
+ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__a211o_1
XANTENNA__09536__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12498__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15979_ net1402 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13635__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13183__A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08520_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[18\] net893
+ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_65_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16647__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17718_ clknet_leaf_81_wb_clk_i _03402_ _01659_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10600__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08451_ net1084 net938 vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__and2_2
XANTENNA__08708__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17649_ clknet_leaf_83_wb_clk_i _03334_ _01590_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08382_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[6\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\]
+ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] _04711_ vssd1 vssd1 vccd1 vccd1
+ _04722_ sky130_fd_sc_hd__nor4_1
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09067__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14060__A2 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18015__1515 vssd1 vssd1 vccd1 vccd1 _18015__1515/HI net1515 sky130_fd_sc_hd__conb_1
XFILLER_0_116_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08814__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_118_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09539__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09003_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[9\] _04799_
+ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11150__B _07489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15838__A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout305_A _07935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1047_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13571__A1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09775__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1214_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 _07795_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16177__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09527__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09905_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[5\] net822 net796 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout512 _05931_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_4
X_17944__1444 vssd1 vssd1 vccd1 vccd1 _17944__1444/HI net1444 sky130_fd_sc_hd__conb_1
Xfanout523 net524 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_2
XANTENNA__17422__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout534 net535 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_2
Xfanout545 _05152_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_2
Xfanout556 net558 vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__buf_2
X_09836_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[13\] net756 net755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__a22o_1
Xfanout567 net568 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_2
Xfanout578 _07753_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_2
Xfanout589 net590 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09571__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout841_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ _06002_ _06036_ _06104_ _06106_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__or4_1
XANTENNA__13626__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17572__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08718_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[5\] net935 vssd1
+ vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__and3_1
XANTENNA__12201__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09698_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[21\] net973 vssd1
+ vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_29_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08502__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08649_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[10\] net906
+ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11660_ net611 _07815_ _07865_ _07864_ vssd1 vssd1 vccd1 vccd1 _07866_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14051__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10611_ net546 _06313_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__nor2_1
X_11591_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\]
+ _07805_ vssd1 vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13330_ net1772 net827 _03806_ _03807_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10542_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] _06881_ net601 vssd1 vssd1
+ vccd1 vccd1 _06882_ sky130_fd_sc_hd__mux2_2
XFILLER_0_122_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15748__A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13261_ _04470_ _03752_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ _05729_ _05736_ vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12212_ net3066 net252 net444 vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__mux2_1
X_15000_ net1179 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__inv_2
X_13192_ net17 net835 net628 net2698 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__o22a_1
XANTENNA_input68_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12143_ net2563 net256 net453 vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__mux2_1
XANTENNA__10915__A3 _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13268__A team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_4__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_88_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09518__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12074_ net2167 net266 net460 vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__mux2_1
X_16951_ clknet_leaf_136_wb_clk_i _02638_ _00934_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09184__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15902_ net1391 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__inv_2
X_11025_ _04948_ net375 vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__nor2_1
X_16882_ clknet_leaf_134_wb_clk_i _02569_ _00865_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12900__A _05654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15833_ net1372 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__inv_2
XANTENNA__13617__A2 _07207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12111__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12825__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10420__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15764_ net1346 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__inv_2
X_12976_ net2914 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[118\] net852 vssd1 vssd1
+ vccd1 vccd1 _02149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17503_ clknet_leaf_24_wb_clk_i _03190_ _01486_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ net1309 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08528__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ net2594 net225 net475 vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__mux2_1
X_15695_ net1213 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11950__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17434_ clknet_leaf_45_wb_clk_i _03121_ _01417_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14646_ net1258 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__inv_2
X_11858_ net1831 net292 net489 vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14042__A2 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08825__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10809_ net525 net519 vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__nor2_1
XANTENNA_19 _07827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17365_ clknet_leaf_124_wb_clk_i _03052_ _01348_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11789_ net2724 net317 net498 vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__mux2_1
X_14577_ net1402 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11251__A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16316_ clknet_leaf_78_wb_clk_i net2983 _00299_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13528_ net198 net194 _07846_ net644 vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17296_ clknet_leaf_15_wb_clk_i _02983_ _01279_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16247_ clknet_leaf_96_wb_clk_i net1796 _00235_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfrtp_1
X_13459_ _03858_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13553__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
X_16178_ clknet_leaf_107_wb_clk_i _01938_ _00166_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__10367__B2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
X_15129_ net1259 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__inv_2
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XANTENNA__09094__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17595__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09391__A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09621_ _05952_ _05953_ _05957_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__or4_2
XANTENNA__13608__A2 _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11619__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[28\] net811 net750 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__a22o_1
XANTENNA__12021__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08503_ net1108 net713 net600 net594 vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_1674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09483_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[30\] net682 _05809_
+ _05811_ _05814_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12956__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout255_A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11860__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08434_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[23\] net919
+ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14033__A2 _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08735__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08365_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\] net764 net621 vssd1
+ vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__o21a_1
XANTENNA__13360__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08454__B net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1164_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ net1134 net971 vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__and2_4
XFILLER_0_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09460__A2 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12691__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1331_A net1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13544__A1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09566__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout791_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08901__C net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout889_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_86_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1307 net1314 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__buf_2
Xfanout320 net321 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1318 net1320 vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_15_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1329 net1341 vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__buf_4
Xfanout331 _06924_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_4
Xfanout342 _06216_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__buf_2
Xfanout353 _03741_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_2
Xfanout364 _03580_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_2
Xfanout375 _06129_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_2
XANTENNA__09920__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 _03570_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09819_ _06158_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__inv_2
Xfanout397 _03567_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_6
XANTENNA__09732__C net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12830_ net1753 net640 net607 _03649_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__a22o_1
X_12761_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[22\] _07154_ net1025 vssd1 vssd1
+ vccd1 vccd1 _03602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1053 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13866__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17318__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11770__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14500_ net1390 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11712_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] _07801_ vssd1 vssd1 vccd1
+ vccd1 _07907_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12692_ net3041 net215 net385 vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__mux2_1
X_15480_ net1178 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14024__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14431_ net1365 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__inv_2
X_11643_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[23\] _07111_ net715 vssd1 vssd1
+ vccd1 vccd1 _07852_ sky130_fd_sc_hd__mux2_1
XANTENNA__12035__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09436__C1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17150_ clknet_leaf_45_wb_clk_i _02837_ _01133_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09987__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16342__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14362_ net1367 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__inv_2
X_11574_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\]
+ vssd1 vssd1 vccd1 vccd1 _07791_ sky130_fd_sc_hd__nor2_2
Xwire710 net711 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10597__A1 _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09179__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09451__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_1
X_16101_ clknet_leaf_92_wb_clk_i _01876_ _00089_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10525_ _06859_ _06860_ _06864_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__or3_1
X_13313_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] net610 _07705_ team_01_WB.instance_to_wrap.cpu.f0.i\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__a31o_1
Xinput39 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
X_17081_ clknet_leaf_51_wb_clk_i _02768_ _01064_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14293_ net1354 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13535__A1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13244_ net3003 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1
+ vccd1 vccd1 _01906_ sky130_fd_sc_hd__a22o_1
X_16032_ clknet_leaf_96_wb_clk_i _01826_ _00026_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10456_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[26\] net741 _06783_ _06784_
+ _06785_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_122_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ net1775 net851 net841 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[1\] vssd1
+ vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a22o_1
X_10387_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[16\] net800 net757 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__a22o_1
XANTENNA__12106__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12126_ net3266 net223 net451 vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17983_ net1483 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__11945__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16934_ clknet_leaf_38_wb_clk_i _02621_ _00917_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12057_ net1988 net293 net463 vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__mux2_1
X_18014__1514 vssd1 vssd1 vccd1 vccd1 _18014__1514/HI net1514 sky130_fd_sc_hd__conb_1
XFILLER_0_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11008_ _05707_ _05932_ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16865_ clknet_leaf_48_wb_clk_i _02552_ _00848_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_15816_ net1311 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__inv_2
X_16796_ clknet_leaf_37_wb_clk_i _02483_ _00779_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15747_ net1187 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__inv_2
X_12959_ net1693 net873 net360 _03714_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10285__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15678_ net1287 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__inv_2
XANTENNA__14015__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13180__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17417_ clknet_leaf_14_wb_clk_i _03104_ _01400_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14629_ net1274 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__inv_2
X_17943__1443 vssd1 vssd1 vccd1 vccd1 _17943__1443/HI net1443 sky130_fd_sc_hd__conb_1
X_08150_ _04604_ _04619_ team_01_WB.instance_to_wrap.cpu.f0.state\[6\] _04516_ vssd1
+ vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__o211a_1
XANTENNA__11234__C1 _05707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17348_ clknet_leaf_52_wb_clk_i _03035_ _01331_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09089__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08081_ _04531_ _04540_ _04545_ _04554_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__or4b_2
XFILLER_0_130_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17279_ clknet_leaf_26_wb_clk_i _02966_ _01262_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16835__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08290__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11537__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12016__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10325__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08983_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[8\] net925 vssd1
+ vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__and3_1
XANTENNA__11855__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09902__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout372_A _06738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08449__B net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[24\] net942
+ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11068__A2 _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09535_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[28\] net978 vssd1
+ vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12686__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1281_A net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_133_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_133_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1379_A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09466_ _05805_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14006__A2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09681__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08417_ net1008 net938 vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__and2_1
XANTENNA__11603__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09397_ _05659_ _05681_ _05707_ _05729_ net560 vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__a41o_1
XFILLER_0_93_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10028__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ net989 net965 vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09433__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1654_A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08279_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] net1683 net1037 vssd1 vssd1
+ vccd1 vccd1 _03408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13517__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10310_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[18\] net802 _06647_
+ _06648_ _06649_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_15_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09296__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11290_ net1155 _04712_ vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__nand2_1
XANTENNA__11528__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10241_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[9\] net814 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__a22o_1
XANTENNA__14930__A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12740__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[10\] net816 net810 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_110_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1104 net1105 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1115 net1116 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__buf_2
XANTENNA__11765__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1126 net1127 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__clkbuf_2
Xfanout1137 net1138 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__clkbuf_2
X_14980_ net1192 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1148 net1149 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__clkbuf_2
Xfanout1159 net1160 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__dlymetal6s2s_1
X_13931_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__and2b_2
Xfanout194 _07634_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17140__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16650_ clknet_leaf_2_wb_clk_i _02337_ _00633_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13862_ net1163 net1058 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[23\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[23\] sky130_fd_sc_hd__and3b_1
XFILLER_0_138_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16708__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15601_ net1293 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12813_ net3125 net640 net607 _03637_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16581_ clknet_leaf_58_wb_clk_i _02268_ _00564_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_104_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12596__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13793_ _04156_ _01833_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15532_ net1219 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[27\] _07566_ net1026 vssd1 vssd1
+ vccd1 vccd1 _03590_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08806__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15463_ net1327 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__inv_2
XANTENNA__13205__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12675_ net2967 net230 net388 vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__mux2_1
XANTENNA__10019__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17202_ clknet_leaf_134_wb_clk_i _02889_ _01185_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14414_ net1338 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__inv_2
X_11626_ net2302 net213 net499 vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__mux2_1
X_15394_ net1266 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09424__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17133_ clknet_leaf_1_wb_clk_i _02820_ _01116_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14345_ net1370 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11557_ net2633 _07787_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13508__A1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire584 _05005_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__buf_4
X_17064_ clknet_leaf_31_wb_clk_i _02751_ _01047_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10508_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[31\] net776 net753 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[31\]
+ _06843_ vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__a221o_1
Xhold609 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11488_ net367 _07771_ net3278 net874 vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__o2bb2a_1
X_14276_ net1367 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09637__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16015_ net1386 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10439_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] net625 _06777_ _06778_
+ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__a22o_2
X_13227_ net2472 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1
+ vccd1 vccd1 _01923_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13158_ net1871 net844 net839 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[18\] vssd1
+ vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16238__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11675__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12109_ net2100 net262 net455 vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__mux2_1
XANTENNA__13456__A _03914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17966_ net1466 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
X_13089_ _03712_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\] net854 vssd1 vssd1
+ vccd1 vccd1 _02036_ sky130_fd_sc_hd__mux2_1
Xhold1309 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16917_ clknet_leaf_123_wb_clk_i _02604_ _00900_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_108_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17897_ net1417 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16848_ clknet_leaf_124_wb_clk_i _02535_ _00831_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17633__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16779_ clknet_leaf_5_wb_clk_i _02466_ _00762_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09320_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[24\] net904
+ net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[24\] vssd1 vssd1 vccd1
+ vccd1 _05660_ sky130_fd_sc_hd__a32o_1
XFILLER_0_34_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08716__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09251_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\] net702 _05585_ _05590_
+ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__o22a_4
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08871__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08202_ net3168 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[71\] net1048 vssd1 vssd1
+ vccd1 vccd1 _03485_ sky130_fd_sc_hd__mux2_1
XANTENNA__17783__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13747__A1 _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09182_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[16\] net660 _05519_
+ _05520_ _05521_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08133_ _04477_ team_01_WB.instance_to_wrap.cpu.f0.num\[17\] team_01_WB.instance_to_wrap.cpu.f0.num\[6\]
+ _04487_ _04594_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__o221a_1
XFILLER_0_126_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout218_A _07835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08064_ _04514_ _04529_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1127_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout587_A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17163__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08966_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[8\] net906 vssd1
+ vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_127_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09282__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[2\] net887 vssd1
+ vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout754_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10497__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09518_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[29\] net803 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[29\]
+ _05846_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__a221o_1
X_10790_ net514 _06957_ _07099_ _07129_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[29\] net701 net656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_135_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12460_ net2579 net218 net413 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__mux2_1
XANTENNA__09406__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18013__1513 vssd1 vssd1 vccd1 vccd1 _18013__1513/HI net1513 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_10_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11411_ _07701_ _07709_ _07728_ net325 vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__o211a_1
XANTENNA__08614__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12391_ net2478 net191 net419 vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14130_ net1685 net604 _04415_ net1169 vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__o211a_1
X_11342_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] net1161 _07670_ vssd1 vssd1 vccd1
+ vccd1 _07671_ sky130_fd_sc_hd__and3_1
XANTENNA__12961__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_112_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14061_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[43\] _04246_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[107\]
+ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__a22o_1
X_11273_ _06100_ _07089_ _06104_ vssd1 vssd1 vccd1 vccd1 _07613_ sky130_fd_sc_hd__a21o_1
XANTENNA__17506__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13012_ net2608 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[82\] net859 vssd1 vssd1
+ vccd1 vccd1 _02113_ sky130_fd_sc_hd__mux2_1
X_10224_ _05264_ _05265_ _05302_ _04750_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__o31a_1
XANTENNA_input50_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17820_ clknet_leaf_66_wb_clk_i net2246 _01760_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09590__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] _06494_ net623 vssd1
+ vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__mux2_1
X_17942__1442 vssd1 vssd1 vccd1 vccd1 _17942__1442/HI net1442 sky130_fd_sc_hd__conb_1
X_17751_ clknet_leaf_64_wb_clk_i _03427_ _01691_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[21\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__16530__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14963_ net1232 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__inv_2
Xhold6 _02018_ vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09192__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10086_ _06422_ _06423_ _06424_ _06425_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__or4_1
XANTENNA__13674__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16702_ clknet_leaf_48_wb_clk_i _02389_ _00685_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13914_ net2996 _04209_ _04210_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_106_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17682_ clknet_leaf_81_wb_clk_i _03366_ _01623_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_14894_ net1284 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16633_ clknet_leaf_46_wb_clk_i _02320_ _00616_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13845_ net1165 net1061 net1773 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[6\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_85_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16680__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16564_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[30\]
+ _00547_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13776_ net1170 _04161_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__nand2_2
X_10988_ net541 _07327_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__or2_1
XANTENNA__09645__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15515_ net1183 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12727_ net1027 _03576_ _03577_ net1161 vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_119_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16495_ clknet_leaf_106_wb_clk_i _02249_ _00478_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14835__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15446_ net1224 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12658_ net2738 net216 net389 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11609_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] _07820_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\]
+ vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__a21o_1
X_15377_ net1291 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12589_ net2871 net192 net397 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17116_ clknet_leaf_37_wb_clk_i _02803_ _01099_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14328_ net1349 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18096_ net637 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_78_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold406 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold417 team_01_WB.instance_to_wrap.a1.ADR_I\[12\] vssd1 vssd1 vccd1 vccd1 net2033
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 net138 vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17186__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17047_ clknet_leaf_140_wb_clk_i _02734_ _01030_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold439 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14259_ net1311 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09664__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout908 _04782_ vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_8
Xfanout919 net921 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_4
X_08820_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[1\] net693 net676 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1106 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1117 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[86\] vssd1 vssd1 vccd1 vccd1
+ net2733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08751_ net1088 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[4\] net913 vssd1
+ vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__and3_1
Xhold1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2744 sky130_fd_sc_hd__dlygate4sd3_1
X_17949_ net1449 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
Xhold1139 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[28\] vssd1 vssd1 vccd1 vccd1
+ net2755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08682_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[7\] net892 vssd1
+ vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__and3_1
XANTENNA__10041__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14090__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08446__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09303_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[22\] net931
+ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12964__S net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11443__A2 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_124_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1077_A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09234_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[21\] net698 net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_131_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08743__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09165_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[16\] net694 net669 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[16\]
+ _05504_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13196__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout502_A _07795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1244_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08116_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] team_01_WB.instance_to_wrap.cpu.f0.num\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__nor2_1
XANTENNA__12943__A2 _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09096_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[13\] net894
+ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__and3_1
XANTENNA__11600__C team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08611__A3 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08047_ net3263 net569 net347 net1064 vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_102_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold940 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[29\] vssd1 vssd1 vccd1 vccd1 net2556
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold951 _02057_ vssd1 vssd1 vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold962 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09574__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold973 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[86\] vssd1 vssd1 vccd1 vccd1
+ net2589 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16553__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold984 _02137_ vssd1 vssd1 vccd1 vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17679__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12204__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] net766 net623 vssd1
+ vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__o21a_1
XANTENNA__10182__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09309__D1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08949_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[6\] net932 vssd1
+ vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_4_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1640 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13120__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3267 sky130_fd_sc_hd__dlygate4sd3_1
X_11960_ net2156 net191 net471 vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__mux2_1
Xhold1662 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[19\] vssd1 vssd1 vccd1 vccd1
+ net3278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1673 team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 net3289
+ sky130_fd_sc_hd__dlygate4sd3_1
X_10911_ _07114_ _07233_ _07239_ _07250_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__a211o_2
XANTENNA__10659__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ net2005 net293 net484 vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__mux2_1
XANTENNA__09740__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11344__A team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13630_ _03883_ _03895_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__nand2_1
X_10842_ _07180_ _07181_ net518 vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__mux2_1
XANTENNA__14081__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17059__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13561_ net980 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _04009_ _04010_
+ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a22o_1
XANTENNA__11434__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08835__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10773_ _06712_ _06740_ _07112_ _06713_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__a31o_1
XANTENNA__14655__A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10642__A0 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15300_ net1239 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__inv_2
X_12512_ net3067 net284 net409 vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16280_ clknet_leaf_76_wb_clk_i _02034_ _00263_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13492_ net712 _04729_ net597 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1
+ vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_97_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15231_ net1254 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__inv_2
XANTENNA__13187__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12443_ net2684 net289 net417 vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08372__B team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12934__A2 _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15162_ net1192 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09260__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12374_ net3161 net231 net424 vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__mux2_1
XANTENNA__10945__A1 _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14113_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[6\] _04265_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__a22o_1
X_11325_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] _07659_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\]
+ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__o21bai_1
X_15093_ net1222 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14044_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[83\] _04251_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11256_ _05681_ net331 _07350_ net369 _07591_ vssd1 vssd1 vccd1 vccd1 _07596_ sky130_fd_sc_hd__o221a_1
X_10207_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[8\] net779 net740 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12114__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ net529 _07237_ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17803_ clknet_leaf_70_wb_clk_i _03479_ _01743_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[73\]
+ sky130_fd_sc_hd__dfrtp_1
X_10138_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[11\] net761 _06476_
+ _06477_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__a211o_1
X_15995_ net1398 vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__inv_2
XANTENNA__11953__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09315__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17734_ clknet_leaf_84_wb_clk_i _03410_ _01674_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_10069_ _06406_ _06408_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14946_ net1262 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__inv_2
XANTENNA__11122__A1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09866__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17665_ clknet_leaf_116_wb_clk_i _03350_ _01606_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14877_ net1250 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16616_ clknet_leaf_24_wb_clk_i _02303_ _00599_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13828_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[21\] net831 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[21\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_63_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17596_ clknet_leaf_69_wb_clk_i _03283_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14072__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09618__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16547_ clknet_leaf_112_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[13\]
+ _00530_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13759_ _04147_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10859__S1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16426__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09659__A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16478_ clknet_leaf_96_wb_clk_i _02232_ _00461_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08563__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15429_ net1209 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__inv_2
XANTENNA__13178__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11189__A1 _06921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16576__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09097__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09397__A4 _05729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold203 team_01_WB.instance_to_wrap.cpu.f0.write_data\[26\] vssd1 vssd1 vccd1 vccd1
+ net1819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold214 team_01_WB.instance_to_wrap.a1.ADR_I\[0\] vssd1 vssd1 vccd1 vccd1 net1830
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold225 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
X_18079_ net1579 vssd1 vssd1 vccd1 vccd1 la_data_out[121] sky130_fd_sc_hd__buf_2
Xhold236 net109 vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[64\] vssd1 vssd1 vccd1 vccd1
+ net1874 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10036__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09921_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[4\] net802 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__a22o_1
Xhold269 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout705 _04758_ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08357__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout716 net717 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__buf_2
XANTENNA__11429__A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ _06188_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__nor2_1
XANTENNA__12024__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout727 net728 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_124_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout738 net739 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10333__A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout749 _04682_ vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__buf_2
X_08803_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[0\] net881 vssd1
+ vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__and3_1
X_09783_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[15\] net787 net783 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__a22o_1
XANTENNA__11863__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18012__1512 vssd1 vssd1 vccd1 vccd1 _18012__1512/HI net1512 sky130_fd_sc_hd__conb_1
X_08734_ _05069_ _05070_ _05073_ net704 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__o32a_2
XFILLER_0_94_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17201__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08665_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[10\] net703 _05001_ _05004_
+ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__o22ai_2
XANTENNA_fanout452_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08457__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1194_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14063__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09609__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08596_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[15\] net698 net697 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[15\]
+ _04922_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12694__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14475__A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout717_A _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10624__B1 _06921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09569__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08473__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16919__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941__1441 vssd1 vssd1 vccd1 vccd1 _17941__1441/HI net1441 sky130_fd_sc_hd__conb_1
XANTENNA__08904__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09217_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[17\] net651 _05532_ _05536_
+ _05538_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12916__A2 _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13574__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08045__A1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[14\] net690 _05459_
+ _05460_ _05475_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_92_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09242__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10927__B2 _06921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08596__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13819__A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09079_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] _04846_ _04845_ vssd1 vssd1
+ vccd1 vccd1 _05419_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11110_ _06404_ _06405_ net345 vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_3__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_12090_ net3063 net291 net460 vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__mux2_1
XANTENNA__09735__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold770 team_01_WB.instance_to_wrap.cpu.f0.num\[29\] vssd1 vssd1 vccd1 vccd1 net2386
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold781 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ _07312_ _07313_ _07380_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold792 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11773__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14800_ net1225 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__inv_2
X_15780_ net1306 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11104__A1 _07064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12992_ net2718 net2688 net852 vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__mux2_1
XANTENNA__09848__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1470 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1481 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[67\] vssd1 vssd1 vccd1 vccd1
+ net3097 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14731_ net1320 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__inv_2
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943_ net2754 net261 net476 vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__mux2_1
XANTENNA__09470__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1492 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net3108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11074__A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17450_ clknet_leaf_2_wb_clk_i _03137_ _01433_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14662_ net1397 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11874_ net1869 net269 net483 vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16401_ clknet_leaf_65_wb_clk_i _02155_ _00384_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[124\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_32_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13613_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\]
+ net597 _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__a31o_1
X_17381_ clknet_leaf_38_wb_clk_i _03068_ _01364_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10825_ _05618_ net331 vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__nor2_1
X_14593_ net1402 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16332_ clknet_leaf_76_wb_clk_i _02086_ _00315_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13544_ net980 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] _03995_ _03996_
+ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09481__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ net336 _07095_ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17844__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16263_ clknet_leaf_107_wb_clk_i net1800 _00251_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11521__B _07784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12109__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13475_ _03929_ _03931_ _03935_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10687_ _06888_ _06892_ net533 vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18002_ net1502 vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_hd__buf_2
XFILLER_0_124_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15214_ net1284 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12426_ net2593 net222 net416 vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09233__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16194_ clknet_leaf_115_wb_clk_i _01954_ _00182_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10918__A1 _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14109__A1 _04348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11948__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15145_ net1228 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13580__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12357_ _07945_ _07946_ net573 vssd1 vssd1 vccd1 vccd1 _07966_ sky130_fd_sc_hd__and3_4
XFILLER_0_121_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10394__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output81_A net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09418__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11308_ net723 _07643_ _07646_ vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__and3_1
X_15076_ net1237 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__inv_2
X_12288_ net2989 net319 net438 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14027_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[10\] _04253_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[114\]
+ _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__a221o_1
XANTENNA__15944__A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11249__A _07588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11239_ _07017_ _07573_ _07578_ _07571_ vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__a211oi_1
XANTENNA__09942__A net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15978_ net1391 vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__inv_2
XANTENNA__09839__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14929_ net1289 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
X_17717_ clknet_leaf_84_wb_clk_i _03401_ _01658_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10600__B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17374__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08450_ net1007 net901 vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__and2_2
XANTENNA__14045__B1 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17648_ clknet_leaf_83_wb_clk_i _03333_ _01589_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08381_ _04624_ _04719_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17579_ clknet_leaf_72_wb_clk_i _03266_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11712__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08814__A3 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12019__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09002_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[9\] net884 vssd1
+ vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11858__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10909__B2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10499__A_N net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13571__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10385__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08232__S net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09904_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[5\] net773 _06241_ _06242_
+ _06243_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__a2111o_1
Xfanout502 _07795_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout513 _05867_ vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__buf_2
Xfanout524 net527 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10137__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout535 net536 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout546 net547 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09852__A _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[13\] net750 net746 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__a22o_1
Xfanout557 net558 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__buf_1
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12689__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout568 _04520_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_4
Xfanout579 net580 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_2
XANTENNA__17717__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _06105_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__inv_2
XANTENNA__08468__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08717_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[5\] net938 vssd1
+ vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__and3_1
XANTENNA__11098__B1 _07339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09290__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09697_ net1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[21\] net966
+ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout834_A team_01_WB.instance_to_wrap.cpu.RU0.next_ihit vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08502__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[10\] net935 vssd1
+ vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14036__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16741__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10937__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08579_ _04885_ _04918_ net600 vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__mux2_2
X_10610_ _06948_ _06949_ net541 vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__mux2_1
X_11590_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _07805_ vssd1 vssd1
+ vccd1 vccd1 _07807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08634__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11341__B _04621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10541_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\] net704 _06870_ _06880_
+ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__o22a_4
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13547__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13260_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] _03751_ vssd1 vssd1 vccd1 vccd1
+ _03752_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10472_ _06811_ vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12211_ net2519 net229 net444 vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__mux2_1
XANTENNA__11768__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13191_ net18 net837 net630 net2198 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ net2418 net259 net452 vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16950_ clknet_leaf_141_wb_clk_i _02637_ _00933_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12073_ net2089 net267 net459 vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11325__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15901_ net1406 vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11024_ net323 _07357_ _07363_ vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__nand3_2
XFILLER_0_99_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16881_ clknet_leaf_15_wb_clk_i _02568_ _00864_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12599__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16271__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13284__A _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15832_ net1372 vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15763_ net1346 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__inv_2
X_12975_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[111\] net2942 net861 vssd1 vssd1
+ vccd1 vccd1 _02150_ sky130_fd_sc_hd__mux2_1
X_17502_ clknet_leaf_46_wb_clk_i _03189_ _01485_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14714_ net1304 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11926_ net2839 net191 net475 vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__mux2_1
XANTENNA__14027__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15694_ net1282 vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ clknet_leaf_47_wb_clk_i _03120_ _01416_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14645_ net1171 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__inv_2
X_11857_ net1735 net314 net490 vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10808_ _07015_ _07099_ _07146_ _07147_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__a211o_1
X_17364_ clknet_leaf_13_wb_clk_i _03051_ _01347_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14576_ net1384 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09454__B1 _04797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11788_ net3103 net319 net498 vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__mux2_1
XANTENNA__13250__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09002__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16315_ clknet_leaf_86_wb_clk_i _02069_ _00298_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[38\]
+ sky130_fd_sc_hd__dfrtp_1
X_13527_ _03942_ _03981_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08662__D1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10739_ _07076_ _07077_ _07078_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__or3b_1
X_17295_ clknet_leaf_143_wb_clk_i _02982_ _01278_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16246_ clknet_leaf_95_wb_clk_i net1770 _00234_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18011__1511 vssd1 vssd1 vccd1 vccd1 _18011__1511/HI net1511 sky130_fd_sc_hd__conb_1
X_13458_ _03914_ _03915_ _03857_ _03859_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11678__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12409_ net2991 net256 net420 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16177_ clknet_leaf_107_wb_clk_i _01937_ _00165_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13389_ _03848_ _03849_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__nor2_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
X_15128_ net1183 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
X_15059_ net1280 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__inv_2
XANTENNA__16614__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10119__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10314__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09672__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08732__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09620_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[24\] net803 net770 _05958_
+ _05959_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a2111o_1
X_17940__1440 vssd1 vssd1 vccd1 vccd1 _17940__1440/HI net1440 sky130_fd_sc_hd__conb_1
XANTENNA__09391__B _05570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10611__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12302__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16764__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08719__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[28\] net758 _05875_ _05879_
+ _05882_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11426__B _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12816__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08502_ net1108 net713 net594 vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10827__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09482_ net1071 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[30\] net900
+ net689 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[30\] vssd1 vssd1 vccd1
+ vccd1 _05822_ sky130_fd_sc_hd__a32o_1
XFILLER_0_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_13__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08433_ net1087 net920 vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__and2_2
XFILLER_0_37_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08735__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ _04693_ _04695_ _04700_ _04703_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__or4_4
XFILLER_0_114_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08227__S net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09445__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13241__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12972__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08295_ net1148 net1151 net1153 net1146 vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__nor4b_2
XANTENNA_fanout415_A _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1157_A team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13529__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16144__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13544__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1324_A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10358__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12752__B1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09285__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16294__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08971__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout310 net312 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_2
Xfanout1308 net1310 vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout321 _07937_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1319 net1320 vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__buf_4
Xfanout332 _06923_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13816__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout354 _03741_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__buf_2
XANTENNA_fanout951_A _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout365 _03580_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__buf_2
Xfanout376 _05262_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_4
X_09818_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] _06157_ net624 vssd1
+ vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__mux2_4
Xfanout387 net390 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_6
XANTENNA__12212__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout398 _03567_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_4
XANTENNA__10521__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09749_ _06085_ _06086_ _06087_ _06088_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__or4_1
XFILLER_0_134_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10818__A0 _07156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12760_ net1825 net639 net606 _03601_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08926__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11711_ net721 _07269_ net615 _07905_ vssd1 vssd1 vccd1 vccd1 _07906_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12691_ net2494 net216 net383 vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14430_ net1361 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__inv_2
X_11642_ net2443 net275 net500 vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__mux2_1
XANTENNA__13232__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_108_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14361_ net1375 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__inv_2
X_11573_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07790_ sky130_fd_sc_hd__nor2_2
XFILLER_0_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11794__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16100_ clknet_leaf_92_wb_clk_i _01875_ _00088_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13312_ net3030 net825 _03791_ _03793_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__o22a_1
XFILLER_0_135_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17080_ clknet_leaf_29_wb_clk_i _02767_ _01063_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10524_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[31\] net682 _06861_
+ _06862_ _06863_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__a2111o_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_1
XFILLER_0_29_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14292_ net1356 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__inv_2
X_16031_ net1362 vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__inv_2
XANTENNA__13279__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13535__A2 _07600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13243_ net3154 net355 net351 net2040 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a22o_1
XANTENNA__16637__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10455_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[26\] net822 net806 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12743__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11546__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13174_ net130 net849 net841 net1811 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10386_ _06723_ _06724_ _06725_ vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__or3_1
XANTENNA__09195__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15494__A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ net3244 net190 net451 vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__mux2_1
X_17982_ net1482 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XANTENNA__13299__A1 _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10134__C net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16787__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16933_ clknet_leaf_40_wb_clk_i _02620_ _00916_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12056_ net2572 net316 net466 vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__mux2_1
XANTENNA__09923__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_9__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _07345_ _07346_ _07344_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12122__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16864_ clknet_leaf_33_wb_clk_i _02551_ _00847_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_15815_ net1311 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__inv_2
X_16795_ clknet_leaf_50_wb_clk_i _02482_ _00778_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11961__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15746_ net1265 vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12958_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[3\] _05219_ net1036 vssd1
+ vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11909_ net3086 net231 net481 vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15677_ net1263 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12889_ _05704_ net578 net362 vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_135_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14628_ net1300 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__inv_2
X_17416_ clknet_leaf_25_wb_clk_i _03103_ _01399_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09427__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13223__B2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17347_ clknet_leaf_18_wb_clk_i _03034_ _01330_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14559_ net1338 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09442__A3 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10309__C net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08080_ _04514_ _04528_ _04532_ _04522_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__o22a_1
XANTENNA__09667__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17278_ clknet_leaf_44_wb_clk_i _02965_ _01261_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16229_ clknet_leaf_105_wb_clk_i net2030 _00217_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10606__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17562__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08290__B net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12734__B1 _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11537__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08953__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08982_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[8\] net906 vssd1
+ vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12032__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10341__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10512__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09603_ net1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[24\] net975
+ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11871__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_A _03580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09534_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[28\] net946 vssd1
+ vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09465_ net601 _05803_ _05804_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_133_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1274_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08416_ net1106 net1109 net1112 net1115 vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__nor4_1
XANTENNA__09418__A0 _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13214__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ _05659_ _05681_ _05707_ net559 vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10028__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08347_ net985 net973 vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__and2_4
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_102_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08481__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08278_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] net1758 net1047 vssd1 vssd1
+ vccd1 vccd1 _03409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout999_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold1647_A team_01_WB.instance_to_wrap.cpu.f0.write_data\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12207__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11528__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10240_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[9\] net749 net739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10171_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[10\] net817 net798 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1105 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1
+ net1105 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1116 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[20\] vssd1 vssd1 vccd1 vccd1
+ net1116 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1127 net1135 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__buf_2
Xfanout1138 net1139 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__clkbuf_2
Xfanout1149 net1150 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13038__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13150__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13930_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__and2b_2
XANTENNA__11347__A team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10251__A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__C1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10503__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout195 net196 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11066__B _06158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13861_ net1163 net1058 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[22\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[22\] sky130_fd_sc_hd__and3b_1
XANTENNA__11466__A1_N net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18010__1510 vssd1 vssd1 vccd1 vccd1 _18010__1510/HI net1510 sky130_fd_sc_hd__conb_1
XFILLER_0_9_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11781__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15600_ net1272 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__inv_2
X_12812_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] net1057 net366 _03636_
+ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__a22o_1
X_16580_ clknet_leaf_54_wb_clk_i _02267_ _00563_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_2_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13792_ _04165_ _04173_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15531_ net1296 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12743_ net2333 net639 net606 _03589_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15462_ net1325 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12674_ net3084 net287 net388 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__mux2_1
XANTENNA__13205__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08880__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08880__B2 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17201_ clknet_leaf_13_wb_clk_i _02888_ _01184_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14413_ net1403 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__inv_2
X_11625_ _07836_ _07837_ net611 vssd1 vssd1 vccd1 vccd1 _07838_ sky130_fd_sc_hd__mux2_2
XANTENNA__15489__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15393_ net1248 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17132_ clknet_leaf_133_wb_clk_i _02819_ _01115_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14344_ net1377 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11556_ team_01_WB.instance_to_wrap.cpu.K0.count\[0\] team_01_WB.instance_to_wrap.cpu.K0.enable
+ _07786_ vssd1 vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08822__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10507_ _06835_ _06844_ _06845_ _06846_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__or4_1
XANTENNA__13508__A2 _07056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17063_ clknet_leaf_123_wb_clk_i _02750_ _01046_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12117__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14275_ net1368 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11487_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[19\] net579 vssd1 vssd1 vccd1
+ vccd1 _07771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16014_ net1373 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09188__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ net2139 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1
+ vccd1 vccd1 _01924_ sky130_fd_sc_hd__a22o_1
X_10438_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\] net764 net621 vssd1
+ vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11956__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13157_ net118 net845 net839 net1619 vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10369_ _04970_ _05379_ _05494_ _05529_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__or4_1
X_12108_ net2838 net231 net457 vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__mux2_1
X_17965_ net1465 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
X_13088_ _03711_ net1717 net858 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__mux2_1
XANTENNA__13141__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15952__A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16916_ clknet_leaf_128_wb_clk_i _02603_ _00899_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12039_ net1981 net235 net464 vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__mux2_1
X_17896_ net1416 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XANTENNA__09950__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16847_ clknet_leaf_143_wb_clk_i _02534_ _00830_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09648__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16778_ clknet_leaf_3_wb_clk_i _02465_ _00761_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15729_ net1324 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_0_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_114_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09250_ _05573_ _05576_ _05587_ _05589_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08201_ net2646 net2881 net1037 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09181_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[16\] net899
+ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10039__C net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12955__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08132_ _04488_ team_01_WB.instance_to_wrap.cpu.f0.num\[5\] _04498_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\]
+ _04595_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_133_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09820__B1 _04749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08063_ _04532_ _04539_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__nor2_1
XANTENNA__12027__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11866__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1022_A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08965_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[8\] net930 vssd1
+ vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout482_A _07949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09563__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13132__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10071__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08896_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[2\] net898 vssd1
+ vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_51_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17458__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12697__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1391_A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout747_A _04682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13382__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09103__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08907__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09517_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[29\] net796 _05844_ _05847_
+ _05849_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13986__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout914_A net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09448_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[29\] net681 net659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[29\]
+ _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13199__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[26\] net701 net666 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__a22o_1
XANTENNA__08923__B net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12946__B1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11410_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] _07693_ vssd1 vssd1 vccd1 vccd1
+ _07728_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_10_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12390_ _07793_ _07946_ net573 vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__and3_1
XANTENNA__09811__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09738__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08642__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11341_ _04511_ _04621_ _07669_ vssd1 vssd1 vccd1 vccd1 _07670_ sky130_fd_sc_hd__and3b_1
XFILLER_0_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14060_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[51\] _04236_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[107\]
+ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11272_ _06100_ _06104_ _07089_ vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__nand3_1
XANTENNA__11776__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ net1976 net1664 net864 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10223_ _06562_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_70_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input43_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\] net767 _06493_ vssd1
+ vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__o21ba_2
XANTENNA__09590__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09473__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13123__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14962_ net1225 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__inv_2
X_17750_ clknet_leaf_56_wb_clk_i _03426_ _01690_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[20\]
+ sky130_fd_sc_hd__dfstp_1
Xhold7 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[8\] vssd1 vssd1 vccd1 vccd1 net1623
+ sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[7\] net794 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__a22o_1
XANTENNA__10412__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16701_ clknet_leaf_49_wb_clk_i _02388_ _00684_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13913_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\] _04209_ net571 vssd1
+ vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_106_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14893_ net1207 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
X_17681_ clknet_leaf_94_wb_clk_i _03365_ _01622_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_134_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13292__A team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16632_ clknet_leaf_28_wb_clk_i _02319_ _00615_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13844_ net1165 net1061 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[5\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[5\] sky130_fd_sc_hd__and3b_1
XANTENNA__12400__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08817__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13775_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\]
+ net604 vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__mux2_1
XANTENNA__13977__A2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16563_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[29\]
+ _00546_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10987_ _06313_ _06339_ net550 vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15514_ net1193 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__inv_2
X_12726_ net1027 team_01_WB.instance_to_wrap.cpu.f0.read_i vssd1 vssd1 vccd1 vccd1
+ _03577_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16494_ clknet_leaf_108_wb_clk_i _02248_ _00477_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16975__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15445_ net1222 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12657_ net2158 net221 net389 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11608_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[30\] _07019_ _04723_ vssd1
+ vssd1 vccd1 vccd1 _07824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15376_ net1271 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08605__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09802__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ _07790_ _07951_ net574 vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__and3_4
XFILLER_0_52_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08552__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17115_ clknet_leaf_48_wb_clk_i _02802_ _01098_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16205__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14327_ net1356 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18095_ net636 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_1
X_11539_ net2952 net1159 net588 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1
+ vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__a22o_1
XANTENNA__10156__A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold407 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[41\] vssd1 vssd1 vccd1 vccd1
+ net2023 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold418 _02010_ vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17046_ clknet_leaf_140_wb_clk_i _02733_ _01029_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold429 _01974_ vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
X_14258_ net1313 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08908__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13209_ net30 net836 net629 net1773 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__o22a_1
XANTENNA__13467__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14189_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[14\] _04457_ vssd1 vssd1 vccd1
+ vccd1 _04458_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout909 net910 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__buf_4
XFILLER_0_81_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09581__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13114__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08750_ net1008 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[4\] net885 vssd1
+ vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__and3_1
Xhold1107 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2723 sky130_fd_sc_hd__dlygate4sd3_1
X_17948_ net1448 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
Xhold1118 team_01_WB.instance_to_wrap.cpu.f0.num\[2\] vssd1 vssd1 vccd1 vccd1 net2734
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13665__A1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_136_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10322__C net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11676__A0 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09333__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08681_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[7\] net882 vssd1
+ vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17879_ clknet_leaf_104_wb_clk_i _03554_ _01819_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08541__B1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12310__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08296__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11428__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_92_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09302_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[22\] net900
+ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[21\] net687 net683 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[21\]
+ _05571_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout230_A _07900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12928__B1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09164_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[16\] net901
+ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08235__S net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08462__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08115_ team_01_WB.instance_to_wrap.cpu.f0.i\[1\] team_01_WB.instance_to_wrap.cpu.f0.num\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12980__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09095_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[13\] net888
+ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17130__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14761__A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1237_A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14145__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_2__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_08046_ net2133 net570 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1
+ vccd1 vccd1 _03545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold930 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold941 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[82\] vssd1 vssd1 vccd1 vccd1
+ net2568 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout697_A _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold963 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10167__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold974 _03492_ vssd1 vssd1 vccd1 vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1404_A net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[10\] vssd1 vssd1 vccd1 vccd1
+ net2612 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09997_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[2\] net752 _06333_ _06334_
+ _06336_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09293__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[6\] net887 vssd1
+ vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_4_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1630 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3246 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09324__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1641 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net3257 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13824__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1652 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[8\] vssd1 vssd1 vccd1 vccd1 net3268
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08879_ _05211_ _05215_ _05218_ net705 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__o32a_4
Xhold1663 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[18\] vssd1 vssd1 vccd1 vccd1
+ net3279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1674 team_01_WB.instance_to_wrap.cpu.f0.state\[8\] vssd1 vssd1 vccd1 vccd1 net3290
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10910_ _07054_ _07235_ _07241_ _07249_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__a31o_1
XANTENNA__12220__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ net2116 net314 net485 vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08637__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ net508 net507 _06636_ _06671_ net548 net537 vssd1 vssd1 vccd1 vccd1 _07181_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11344__B team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13560_ net722 _07171_ net1066 vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10772_ _06598_ _06604_ _06742_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__a21o_1
XANTENNA__08934__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17909__1601 vssd1 vssd1 vccd1 vccd1 net1601 _17909__1601/LO sky130_fd_sc_hd__conb_1
XFILLER_0_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12511_ net2588 net251 net408 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10642__A1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16228__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13491_ _03841_ _03842_ _03950_ _03839_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15230_ net1248 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__inv_2
X_12442_ net2843 net257 net417 vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15161_ net1305 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12373_ net2634 net264 net425 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__mux2_1
XANTENNA__12890__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14112_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[38\] _04230_ _04259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__a22o_1
XANTENNA__10945__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16378__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14136__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09765__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11324_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\]
+ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] _07658_ vssd1 vssd1 vccd1 vccd1
+ _07659_ sky130_fd_sc_hd__or4_1
X_15092_ net1291 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17623__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14043_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] _04249_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[115\]
+ _04331_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11255_ net523 _07534_ _07594_ vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10158__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[8\] net949 vssd1
+ vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11519__B net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11186_ _07234_ _07483_ net525 vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17802_ clknet_leaf_85_wb_clk_i net2882 _01742_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_10137_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[11\] net810 net782 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__a22o_1
XANTENNA__13647__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15994_ net1391 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09315__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17733_ clknet_leaf_81_wb_clk_i _03409_ _01673_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11658__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10068_ _06285_ _06407_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14945_ net1243 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12130__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17664_ clknet_leaf_116_wb_clk_i _03349_ _01605_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_82_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14876_ net1174 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09005__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16615_ clknet_leaf_16_wb_clk_i _02302_ _00598_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08547__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13827_ net2160 net831 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[20\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09079__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17595_ clknet_leaf_69_wb_clk_i _03282_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13758_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 _04147_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_128_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16546_ clknet_leaf_110_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[12\]
+ _00529_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ net3133 net251 net384 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17153__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13689_ team_01_WB.instance_to_wrap.cpu.c0.count\[6\] team_01_WB.instance_to_wrap.cpu.c0.count\[5\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[15\] team_01_WB.instance_to_wrap.cpu.c0.count\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__or4bb_1
X_16477_ clknet_leaf_95_wb_clk_i _02231_ _00460_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15428_ net1237 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15359_ net1256 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09251__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold204 net110 vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09675__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14127__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold215 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
X_18078_ net1578 vssd1 vssd1 vccd1 vccd1 la_data_out[120] sky130_fd_sc_hd__buf_2
Xhold226 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 _01976_ vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09920_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[4\] net807 net772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__a22o_1
Xhold248 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ clknet_leaf_39_wb_clk_i _02716_ _01012_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold259 _02103_ vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09394__B _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10149__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12305__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10614__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout706 net709 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_6
XFILLER_0_111_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09851_ _05454_ _06190_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__xnor2_1
Xfanout717 _04723_ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_2
XANTENNA__09554__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout728 net729 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_124_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 _04686_ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_6
X_08802_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[0\] net879 vssd1
+ vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__and3_1
X_09782_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[15\] net820 _06120_
+ _06121_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13638__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08733_ _05061_ _05064_ _05071_ _05072_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__or4_1
XANTENNA__09306__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08664_ _04995_ _04996_ _05002_ _05003_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__or4_1
XANTENNA__12040__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _04932_ _04933_ _04934_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_137_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout445_A _07959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1187_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout612_A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08473__B net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1354_A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09216_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[17\] net655 _05535_
+ _05542_ _05553_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16520__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09288__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09147_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[14\] net682 _05467_
+ _05472_ net709 vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_92_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09242__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10388__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14118__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13819__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] _04846_ _04845_ vssd1 vssd1
+ vccd1 vccd1 _05418_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout981_A _04499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08029_ team_01_WB.instance_to_wrap.cpu.f0.state\[7\] net569 vssd1 vssd1 vccd1 vccd1
+ _04525_ sky130_fd_sc_hd__nor2_2
XANTENNA__16670__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12215__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17796__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold760 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[40\] vssd1 vssd1 vccd1 vccd1
+ net2376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 team_01_WB.instance_to_wrap.cpu.f0.write_data\[12\] vssd1 vssd1 vccd1 vccd1
+ net2398 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ _07295_ _07296_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__nor2_1
XANTENNA__09545__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold793 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[42\] vssd1 vssd1 vccd1 vccd1
+ net2409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11339__B _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13629__A1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12991_ net1805 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[103\] net862 vssd1 vssd1
+ vccd1 vccd1 _02134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11104__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13046__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1460 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 net3076
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08505__B1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1471 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14730_ net1351 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11942_ net3212 net233 net477 vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10312__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1482 team_01_WB.instance_to_wrap.cpu.c0.count\[11\] vssd1 vssd1 vccd1 vccd1 net3098
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1493 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3109 sky130_fd_sc_hd__dlygate4sd3_1
X_14661_ net1382 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__inv_2
XANTENNA__10863__B2 _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11873_ net2249 net237 net483 vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__mux2_1
X_16400_ clknet_leaf_72_wb_clk_i net1912 _00383_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_13612_ _03888_ _04052_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10824_ _05619_ net507 vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__nand2_1
X_14592_ net1384 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__inv_2
X_17380_ clknet_leaf_51_wb_clk_i _03067_ _01363_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10615__A1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16331_ clknet_leaf_75_wb_clk_i net2466 _00314_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13543_ net722 _07111_ net1066 vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10755_ _04844_ net510 vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16262_ clknet_leaf_105_wb_clk_i _02022_ _00250_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10091__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13474_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _05592_ _05616_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__a22o_1
X_10686_ _06979_ _07025_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_1419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09198__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18001_ net1501 vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_hd__buf_2
X_15213_ net1212 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12425_ net3022 net223 net415 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16193_ clknet_leaf_115_wb_clk_i _01953_ _00181_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10379__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14109__A2 _04395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15144_ net1276 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12356_ net2284 net291 net428 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09784__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08830__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11307_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _05116_ vssd1 vssd1 vccd1
+ vccd1 _07646_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15075_ net1186 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12287_ net2319 net308 net438 vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__mux2_1
XANTENNA__12125__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14026_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[98\] _04244_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[58\]
+ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__a22o_1
X_11238_ net553 _07266_ _07572_ _07575_ _07577_ vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09536__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11964__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10551__A0 _06707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ _07269_ _07290_ _07308_ _07508_ vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_93_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10570__A_N _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15977_ net1339 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17716_ clknet_leaf_84_wb_clk_i _03400_ _01657_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17519__CLK clknet_leaf_143_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14928_ net1225 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
X_18085__1585 vssd1 vssd1 vccd1 vccd1 _18085__1585/HI net1585 sky130_fd_sc_hd__conb_1
XFILLER_0_117_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10303__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17647_ clknet_leaf_83_wb_clk_i _03332_ _01588_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14859_ net1295 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08380_ _04624_ _04719_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17578_ clknet_leaf_77_wb_clk_i _03265_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17669__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16529_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[27\]
+ _00512_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17887__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10082__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09001_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[9\] net903 vssd1
+ vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09224__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09775__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08740__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13308__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12035__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10344__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17049__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09903_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[5\] net815 net745 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_6_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout503 _06857_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__clkbuf_4
Xfanout514 net515 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_4
Xfanout525 net526 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17908__1600 vssd1 vssd1 vccd1 vccd1 net1600 _17908__1600/LO sky130_fd_sc_hd__conb_1
Xfanout536 _05190_ vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout395_A _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11874__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout547 _05152_ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_2
X_09834_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[13\] net800 net768 vssd1
+ vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_127_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10542__A0 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1102_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout558 _05114_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08749__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10998__B _05263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout569 net570 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09765_ net507 _06099_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09571__C net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout562_A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__B net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[5\] net928 vssd1
+ vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__and3_1
X_09696_ _06034_ _06035_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[10\] net885
+ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14486__A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13390__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08578_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] net702 _04900_ _04917_
+ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__o22a_4
XANTENNA__08484__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09463__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10540_ _06875_ _06877_ _06878_ _06879_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__or4_1
XFILLER_0_119_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10471_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] net625 _06809_ _06810_
+ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__a22o_4
XANTENNA__10443__A_N net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15110__A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12210_ net2166 net288 net446 vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13190_ net19 net835 net628 net1984 vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08650__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12770__A1 _07135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ net2818 net231 net452 vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__mux2_1
XANTENNA__10254__A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09518__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12072_ net2271 net238 net459 vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold590 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11784__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15900_ net1388 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__inv_2
XANTENNA__16416__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11023_ _07361_ _07362_ _07223_ _07359_ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__a211oi_1
X_16880_ clknet_leaf_128_wb_clk_i _02567_ _00863_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10533__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15831_ net1372 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12974_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[112\] net1832 net860 vssd1 vssd1
+ vccd1 vccd1 _02151_ sky130_fd_sc_hd__mux2_1
X_15762_ net1321 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09151__A0 _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12825__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10420__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16566__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17501_ clknet_leaf_49_wb_clk_i _03188_ _01484_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1290 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14713_ net1304 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__inv_2
X_11925_ _07790_ net576 _07946_ vssd1 vssd1 vccd1 vccd1 _07950_ sky130_fd_sc_hd__and3_1
X_15693_ net1208 vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17432_ clknet_leaf_29_wb_clk_i _03119_ _01415_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ net2653 net318 net490 vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__mux2_1
X_14644_ net1196 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08825__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ _07004_ _07100_ net329 _06988_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__a22o_1
X_14575_ net1339 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__inv_2
X_17363_ clknet_leaf_137_wb_clk_i _03050_ _01346_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11787_ net2211 net307 net498 vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16314_ clknet_leaf_61_wb_clk_i _02068_ _00297_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[37\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10738_ _06964_ _07055_ _07068_ net530 vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13526_ _03851_ _03852_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__nand2_1
X_17294_ clknet_leaf_6_wb_clk_i _02981_ _01277_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13457_ _03859_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__or2_1
X_16245_ clknet_leaf_95_wb_clk_i net1729 _00233_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
X_10669_ _07006_ _07008_ net541 vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12408_ net2525 net262 net421 vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16176_ clknet_leaf_107_wb_clk_i _01936_ _00164_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13388_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _05727_ vssd1 vssd1
+ vccd1 vccd1 _03849_ sky130_fd_sc_hd__nor2_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_50_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XANTENNA__12761__A1 _07154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
X_15127_ net1195 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__inv_2
X_12339_ net3108 net269 net427 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__mux2_1
XANTENNA__10164__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15058_ net1234 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__inv_2
XANTENNA__11694__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14009_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[121\] _04250_ _04297_ _04299_
+ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__a211o_1
XANTENNA__17341__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09390__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16909__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10611__B _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09550_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[28\] net794 _05873_ _05877_
+ _05878_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_95_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08501_ net730 _04752_ _04838_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1
+ vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__o31a_1
XANTENNA__10827__A1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09481_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[30\] net698 net697 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08432_ net1007 net925 vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__and2_2
XFILLER_0_56_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08363_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[30\] net739 _04701_
+ _04702_ net768 vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09445__A1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09996__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ net1127 net973 vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__and2_4
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11869__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1052_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09748__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09566__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12752__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10074__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_2
Xfanout311 net312 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_1
XFILLER_0_111_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout777_A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1309 net1310 vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__buf_4
XFILLER_0_10_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout333 _06923_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_2
Xfanout344 _04748_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08479__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout355 net356 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16589__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout366 _03580_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09381__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09817_ _06149_ _06153_ _06155_ _06156_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__o31a_4
XANTENNA__09920__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout377 _04969_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_4
Xfanout388 net389 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_6
XFILLER_0_96_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout944_A _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout399 _03566_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_6
XFILLER_0_119_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09748_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[20\] net803 _06070_
+ _06078_ _06080_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_97_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13832__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09679_ _06016_ _06017_ _06018_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08487__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11710_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[9\] net717 vssd1 vssd1 vccd1
+ vccd1 _07905_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_95_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08926__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12690_ net2584 net220 net385 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08645__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11641_ _07848_ _07849_ _07850_ net611 vssd1 vssd1 vccd1 vccd1 _07851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10046__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14360_ net1375 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__inv_2
XANTENNA__09987__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11572_ _04726_ _04752_ _04846_ vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__or3_2
XFILLER_0_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11779__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13311_ net565 _07709_ _03792_ net829 vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__a31o_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_10523_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[31\] net926 vssd1
+ vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14291_ net1382 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16030_ net1362 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__inv_2
X_13242_ net2739 net355 net351 net1064 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a22o_1
X_10454_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[26\] net976
+ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__and3_1
XANTENNA_input73_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18084__1584 vssd1 vssd1 vccd1 vccd1 _18084__1584/HI net1584 sky130_fd_sc_hd__conb_1
XFILLER_0_66_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12743__B2 _03589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13173_ net133 net850 net842 net1693 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10385_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[16\] net761 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__a22o_1
XANTENNA__17364__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10415__C net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12124_ _07791_ net575 _07793_ vssd1 vssd1 vccd1 vccd1 _07957_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17981_ net1481 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_44_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12055_ net2103 net318 net466 vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__mux2_1
X_16932_ clknet_leaf_51_wb_clk_i _02619_ _00915_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12403__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09372__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ _05729_ _06812_ vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16863_ clknet_leaf_8_wb_clk_i _02550_ _00846_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_15814_ net1311 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__inv_2
X_16794_ clknet_leaf_45_wb_clk_i _02481_ _00777_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15745_ net1249 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__inv_2
X_12957_ net1751 net872 net359 _03713_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15015__A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_104_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11908_ net2273 net264 net481 vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10285__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15676_ net1174 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12888_ net1857 net870 net357 _03666_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09013__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17415_ clknet_leaf_123_wb_clk_i _03102_ _01398_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14627_ net1295 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11839_ net2162 net242 net487 vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14854__A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11234__A1 _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17346_ clknet_leaf_36_wb_clk_i _03033_ _01329_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09948__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14558_ net1336 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08852__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11689__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13509_ _03966_ _03967_ net1067 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_43_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17277_ clknet_leaf_40_wb_clk_i _02964_ _01260_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14489_ net1399 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16228_ clknet_leaf_107_wb_clk_i net1708 _00216_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10606__B _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11537__A2 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12734__B2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16159_ clknet_leaf_98_wb_clk_i _01922_ _00147_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10745__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10325__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08981_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[8\] net902 vssd1
+ vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__and3_1
XANTENNA__10840__S0 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16731__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12313__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08299__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09902__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_143_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09602_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[24\] net974
+ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__and3_1
XANTENNA__16881__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09533_ net1126 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[28\] net976
+ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout358_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ net599 _05802_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__or2_1
XANTENNA__10276__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08465__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08415_ net712 _04751_ _04752_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__or3_4
XFILLER_0_93_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09395_ _05659_ _05681_ net559 vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1267_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10028__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ net1129 net941 vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08277_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\] net3006 net1037 vssd1 vssd1
+ vccd1 vccd1 _03410_ sky130_fd_sc_hd__mux2_1
XANTENNA__16261__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17387__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08481__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09296__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout894_A _04793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11528__A2 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_142_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_142_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09593__A _05707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10170_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[10\] net805 net769 vssd1
+ vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_110_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13827__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11628__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1106 net1107 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__buf_2
Xfanout1117 net1118 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__clkbuf_2
Xfanout1128 net1129 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__buf_2
Xfanout1139 net1142 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__buf_2
XANTENNA__09354__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08002__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout185 net186 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout196 _07634_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11757__A_N team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13860_ net1163 net1058 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[21\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[21\] sky130_fd_sc_hd__and3b_1
XFILLER_0_57_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08937__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13989__B1 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[6\] _07323_ net1033 vssd1 vssd1
+ vccd1 vccd1 _03636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13791_ _01834_ _01833_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11363__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ net1273 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12742_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] net1054 net363 _03588_
+ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12673_ net2990 net255 net387 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__mux2_1
X_15461_ net1207 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__inv_2
XANTENNA__13205__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16604__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17200_ clknet_leaf_127_wb_clk_i _02887_ _01183_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10019__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14412_ net1403 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__inv_2
X_11624_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _07819_ vssd1 vssd1
+ vccd1 vccd1 _07837_ sky130_fd_sc_hd__xor2_1
X_15392_ net1242 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08672__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12964__A1 _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17131_ clknet_leaf_0_wb_clk_i _02818_ _01114_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11555_ net1168 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.next_state
+ sky130_fd_sc_hd__inv_2
XFILLER_0_52_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14343_ net1373 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10506_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[31\] net815 net805 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__a22o_1
X_17062_ clknet_leaf_42_wb_clk_i _02749_ _01045_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14274_ net1368 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11486_ net367 _07770_ net2111 net874 vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__16754__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16013_ net1385 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13225_ net3059 net355 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1
+ vccd1 vccd1 _01925_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10437_ _06766_ _06768_ _06773_ _06776_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__or4_2
XFILLER_0_46_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ net120 net845 net839 net2308 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10368_ _06707_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12107_ net2201 net263 net456 vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__mux2_1
X_17964_ net1464 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
XANTENNA__12133__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10442__A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13087_ _03710_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\] net863 vssd1 vssd1
+ vccd1 vccd1 _02038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10299_ net505 _06638_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__nand2_1
XANTENNA__13141__A1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09008__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16915_ clknet_leaf_135_wb_clk_i _02602_ _00898_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12038_ net2449 net242 net464 vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__mux2_1
X_17895_ net1598 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XANTENNA__11972__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16846_ clknet_leaf_5_wb_clk_i _02533_ _00829_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16134__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16777_ clknet_leaf_9_wb_clk_i _02464_ _00760_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13989_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[72\] _04235_ _04254_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[96\]
+ _04271_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15728_ net1223 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15659_ net1298 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__inv_2
XANTENNA__16284__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08871__A2 _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08200_ net1629 net2227 net1050 vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11207__A1 _06915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11207__B2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09180_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[16\] net888
+ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13601__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08582__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08131_ _04465_ team_01_WB.instance_to_wrap.cpu.f0.num\[31\] team_01_WB.instance_to_wrap.cpu.f0.num\[26\]
+ _04469_ _04588_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17329_ clknet_leaf_15_wb_clk_i _03016_ _01312_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11720__B _07308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12308__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09820__A1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08623__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08062_ _04513_ team_01_WB.instance_to_wrap.cpu.K0.code\[1\] team_01_WB.instance_to_wrap.cpu.K0.code\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__or3b_2
XFILLER_0_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10430__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_1__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12043__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[8\] net892 vssd1
+ vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1015_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08139__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09336__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08895_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[2\] net903 vssd1
+ vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_51_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11882__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11694__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10497__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08757__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12891__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1384_A net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16627__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18083__1583 vssd1 vssd1 vccd1 vccd1 _18083__1583/HI net1583 sky130_fd_sc_hd__conb_1
XANTENNA__10249__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09516_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[29\] net813 net770 _05840_
+ _05843_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11446__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[29\] net673 net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a22o_1
XANTENNA__14494__A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout907_A net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09378_ _05716_ _05717_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12946__A1 _05337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08329_ net989 net951 vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12218__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10957__A0 _06912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08614__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09272__C1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14148__B1 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11340_ _07651_ team_01_WB.instance_to_wrap.cpu.f0.state\[6\] _04576_ vssd1 vssd1
+ vccd1 vccd1 _07669_ sky130_fd_sc_hd__or3b_1
XFILLER_0_6_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11271_ _07601_ _07602_ _07610_ vssd1 vssd1 vccd1 vccd1 _07611_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13010_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[76\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[84\]
+ net856 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__mux2_1
X_10222_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] net627 _06560_ _06561_
+ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__a22o_2
XANTENNA__09575__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10153_ _06486_ _06490_ _06492_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__nor3_1
XANTENNA__09327__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14961_ net1289 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__inv_2
XANTENNA_input36_A gpio_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[7\] net791 net747 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_1594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11792__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[25\] vssd1 vssd1 vccd1 vccd1 net1624
+ sky130_fd_sc_hd__dlygate4sd3_1
X_16700_ clknet_leaf_37_wb_clk_i _02387_ _00683_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_58_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13912_ _04209_ net571 _04208_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_106_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17680_ clknet_leaf_94_wb_clk_i _03364_ _01621_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_106_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14892_ net1205 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16631_ clknet_leaf_138_wb_clk_i _02318_ _00614_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13843_ net1165 net1060 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[4\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[4\] sky130_fd_sc_hd__and3b_1
XFILLER_0_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11093__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17552__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16562_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[28\]
+ _00545_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13774_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ _04146_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__mux2_1
X_10986_ _07012_ _07325_ net541 vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15513_ net1260 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__inv_2
X_12725_ team_01_WB.instance_to_wrap.cpu.DM0.state\[0\] _07783_ team_01_WB.instance_to_wrap.cpu.DM0.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16493_ clknet_leaf_106_wb_clk_i _02247_ _00476_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12917__A _05564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09498__A _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15444_ net1288 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__inv_2
X_12656_ net3045 net224 net387 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08833__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11607_ net2841 net192 net499 vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15375_ net1213 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__inv_2
X_12587_ net2124 net292 net400 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12128__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08605__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17114_ clknet_leaf_60_wb_clk_i _02801_ _01097_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14139__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14326_ net1358 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11538_ net2255 net1159 net589 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] vssd1
+ vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__a22o_1
X_18094_ net636 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold408 _03455_ vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11967__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17045_ clknet_leaf_125_wb_clk_i _02732_ _01028_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold419 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[28\] net580 vssd1 vssd1 vccd1
+ vccd1 _07762_ sky130_fd_sc_hd__nand2_1
X_14257_ net1313 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13208_ net31 net836 net629 net2850 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14188_ net1410 _04456_ _04457_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__nor3_1
XANTENNA__09664__C net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13139_ net1767 net850 net632 team_01_WB.instance_to_wrap.a1.ADR_I\[4\] vssd1 vssd1
+ vccd1 vccd1 _02002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1108 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2724 sky130_fd_sc_hd__dlygate4sd3_1
X_17947_ net1447 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
Xhold1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2735 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13665__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11676__A1 _07541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08680_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[7\] net923 vssd1
+ vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__and3_1
X_17878_ clknet_leaf_109_wb_clk_i _03553_ _01818_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08541__B2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16829_ clknet_leaf_40_wb_clk_i _02516_ _00812_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08296__B net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14090__A2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09301_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[22\] net900 vssd1
+ vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08844__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09232_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[21\] net691 net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08743__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12928__A1 _05490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09201__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09163_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[16\] net655 _05500_
+ _05501_ _05502_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08057__B1 _04534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12038__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10347__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08114_ team_01_WB.instance_to_wrap.cpu.f0.i\[11\] team_01_WB.instance_to_wrap.cpu.f0.num\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09094_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[13\] net914 vssd1
+ vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11877__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08045_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[10\] net569 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__a22o_1
Xhold920 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[119\] vssd1 vssd1 vccd1 vccd1
+ net2536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold931 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1132_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold942 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09557__B1 _05896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold953 _03488_ vssd1 vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13353__B2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold964 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09574__C net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17425__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold975 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1
+ net2602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08765__D1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15873__A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold997 _02041_ vssd1 vssd1 vccd1 vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09996_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[2\] net763 _06317_ _06335_
+ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08947_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[6\] net939 vssd1
+ vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__and3_1
XANTENNA__14489__A net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1620 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3236 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1631 team_01_WB.instance_to_wrap.a1.ADR_I\[2\] vssd1 vssd1 vccd1 vccd1 net3247
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11667__A1 _07251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10810__A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12501__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1642 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1653 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3269 sky130_fd_sc_hd__dlygate4sd3_1
X_08878_ _05208_ _05212_ _05216_ _05217_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__or4_1
Xhold1664 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 net3280
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1675 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 net3291
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10840_ net375 _06158_ _06707_ net372 net549 net533 vssd1 vssd1 vccd1 vccd1 _07180_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_131_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14081__A2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13840__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ net562 _07092_ _07093_ _07110_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__a31o_2
XANTENNA__08835__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12510_ net2949 net229 net408 vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13490_ _03842_ _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_118_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12441_ net2921 net260 net418 vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__mux2_1
XANTENNA__08653__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08048__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09796__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13592__A1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15160_ net1172 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12372_ net2752 net267 net423 vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09260__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11787__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14111_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[102\] _04244_ _04247_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[70\]
+ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__a22o_1
XANTENNA__10945__A3 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11323_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\]
+ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\] team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\]
+ vssd1 vssd1 vccd1 vccd1 _07658_ sky130_fd_sc_hd__or4_1
X_15091_ net1280 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14042_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\] _04265_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[27\]
+ _04330_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__a221o_1
X_11254_ _06906_ _07081_ _07084_ _05263_ net339 vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__o221a_1
XFILLER_0_43_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08161__S net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10158__A1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10704__B net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[8\] net962 vssd1
+ vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11185_ _07375_ _07523_ _07524_ net339 vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17801_ clknet_leaf_77_wb_clk_i net3251 _01741_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_10136_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[11\] net820 net804 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__a22o_1
X_15993_ net1338 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13647__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17732_ clknet_leaf_84_wb_clk_i _03408_ _01672_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10067_ _06280_ _06283_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__or2_1
X_14944_ net1241 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__inv_2
XANTENNA__11658__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12411__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08828__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09720__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17663_ clknet_leaf_114_wb_clk_i _03348_ _01604_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16942__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10330__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14875_ net1184 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16614_ clknet_leaf_39_wb_clk_i _02301_ _00597_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_82_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13826_ net2551 net831 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[19\]
+ sky130_fd_sc_hd__and2_1
X_17594_ clknet_leaf_69_wb_clk_i _03281_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10881__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14072__A2 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16545_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[11\]
+ _00528_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13757_ _04141_ _04142_ _04145_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__and3_2
XANTENNA__13846__A_N net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13280__B1 _04621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10969_ _06255_ _06410_ _07291_ vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_75_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10094__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12708_ net2913 net229 net384 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16476_ clknet_leaf_95_wb_clk_i _02230_ _00459_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13688_ team_01_WB.instance_to_wrap.cpu.c0.count\[15\] _04109_ vssd1 vssd1 vccd1
+ vccd1 _04111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08563__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15427_ net1188 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__inv_2
XANTENNA__08039__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12639_ net2195 net259 net393 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13583__A1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16322__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15358_ net1271 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17448__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08860__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09251__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold205 _01977_ vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
X_14309_ net1350 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18077_ net1577 vssd1 vssd1 vccd1 vccd1 la_data_out[119] sky130_fd_sc_hd__buf_2
XFILLER_0_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold216 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[120\] vssd1 vssd1 vccd1 vccd1
+ net1832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15289_ net1260 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold227 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold238 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[20\] vssd1 vssd1 vccd1 vccd1
+ net1854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17028_ clknet_leaf_51_wb_clk_i _02715_ _01011_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold249 team_01_WB.instance_to_wrap.a1.ADR_I\[18\] vssd1 vssd1 vccd1 vccd1 net1865
+ sky130_fd_sc_hd__dlygate4sd3_1
X_18082__1582 vssd1 vssd1 vccd1 vccd1 _18082__1582/HI net1582 sky130_fd_sc_hd__conb_1
XFILLER_0_81_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_84_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17598__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ net377 _05378_ _05416_ net561 vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__a31o_1
Xfanout707 net709 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_8
Xfanout718 net719 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_124_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout729 _04720_ vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_124_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[0\] net913 vssd1
+ vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__and3_1
X_09781_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[15\] net738 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12321__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08732_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[5\] net664 _05048_ _05050_
+ _05055_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_98_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10630__A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09711__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08738__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[10\] net657 _04982_
+ _04984_ _04992_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_94_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08594_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[15\] net904
+ net693 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[15\] vssd1 vssd1 vccd1
+ vccd1 _04934_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_137_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14063__A2 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_93_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08278__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1082_A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16029__A net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout438_A _07963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10085__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09490__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09569__C net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09215_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[17\] net685 _05534_
+ _05537_ _05550_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_49_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10077__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout605_A _04151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1347_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ _05482_ _05483_ _05484_ _05485_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__or4_2
XANTENNA__13574__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13388__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09077_ _05416_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16815__CLK clknet_leaf_143_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08028_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid _04523_ vssd1 vssd1 vccd1 vccd1
+ _04524_ sky130_fd_sc_hd__nand2_4
Xhold750 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[26\] vssd1 vssd1 vccd1 vccd1
+ net2366 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout974_A _04633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold761 _02079_ vssd1 vssd1 vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[0\] vssd1 vssd1 vccd1 vccd1 net2410
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16965__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[2\] net787 net780 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13629__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12231__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ net2736 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[104\] net860 vssd1 vssd1
+ vccd1 vccd1 _02135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1450 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3066 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08648__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1461 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3077 sky130_fd_sc_hd__dlygate4sd3_1
X_11941_ net2339 net265 net476 vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__mux2_1
Xhold1472 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[31\] vssd1 vssd1 vccd1 vccd1
+ net3088 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14039__C1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1483 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3099 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13869__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1494 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net3110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14660_ net1382 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11872_ net2340 net241 net483 vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13611_ _03897_ _04051_ _03891_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__a21oi_1
X_10823_ _07055_ _07161_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__nor2_1
X_14591_ net1339 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08808__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16330_ clknet_leaf_61_wb_clk_i _02084_ _00313_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[53\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_113_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13542_ net185 _03993_ _03994_ net725 vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_1346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10754_ _04844_ _05996_ vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__or2_1
XANTENNA__09481__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16261_ clknet_leaf_107_wb_clk_i net1826 _00249_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
X_10685_ net515 _07023_ _07024_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__and3_1
X_13473_ _03855_ _03921_ _03933_ _03853_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18000_ net1500 vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_hd__buf_2
XANTENNA__10418__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13565__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09769__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15212_ net1182 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__inv_2
X_12424_ net3132 net189 net415 vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__mux2_1
X_16192_ clknet_leaf_115_wb_clk_i _01952_ _00180_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09233__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15143_ net1327 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16495__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13298__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ net2322 net316 net430 vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__mux2_1
XANTENNA__12406__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10715__A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11306_ _07645_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] _07638_ vssd1
+ vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12286_ net2144 net309 net436 vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15074_ net1268 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14025_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[10\] _04226_ _04251_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[82\]
+ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__a221o_1
X_11237_ net523 _07219_ _07576_ vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__o21a_1
X_11168_ _07323_ _07438_ _07491_ _07507_ vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_8_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10551__A1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10119_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[6\] net806 net759 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12141__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15976_ net1336 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__inv_2
X_11099_ _06406_ _06408_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__and2_1
XANTENNA__12828__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09016__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17715_ clknet_leaf_84_wb_clk_i _03399_ _01656_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08558__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14927_ net1212 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
XANTENNA__11980__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17120__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17646_ clknet_leaf_83_wb_clk_i _03331_ _01587_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14858_ net1282 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14045__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08855__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12056__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13809_ net3128 net833 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[2\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_54_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17577_ clknet_leaf_72_wb_clk_i _03264_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10596__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14789_ net1205 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16528_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[26\]
+ _00511_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11803__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17270__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16459_ clknet_leaf_6_wb_clk_i _02213_ _00442_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09000_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[9\] net932 vssd1
+ vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__and3_1
XANTENNA__16838__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09224__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12316__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13308__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[5\] net789 net776 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_1662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout504 _06779_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__buf_2
Xfanout515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout526 net527 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_2
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09833_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[13\] net821 net794 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__a22o_1
Xfanout537 net538 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_4
Xfanout548 net549 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout290_A _07896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10542__A1 _06881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout559 net561 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16218__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10998__C _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12051__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ _06068_ _06069_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08715_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[5\] net932 vssd1
+ vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__and3_1
XANTENNA__13492__B1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09695_ net509 _06033_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__nor2_1
XANTENNA__11890__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1297_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08646_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[10\] net909
+ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14036__A2 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08577_ _04904_ _04908_ _04912_ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout722_A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10058__B1 _06396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09299__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09463__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13547__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09596__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10470_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\] net764 net621 vssd1
+ vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__o21a_1
XANTENNA__09215__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08931__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09129_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[14\] net880
+ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__and3_1
XANTENNA__12226__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12140_ net2857 net264 net453 vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12071_ net2056 net239 net459 vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__mux2_1
Xhold580 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold591 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _05529_ net372 vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11366__A team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15830_ net1372 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10270__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15761_ net1321 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__inv_2
X_12973_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[113\] net1913 net866 vssd1 vssd1
+ vccd1 vccd1 _02152_ sky130_fd_sc_hd__mux2_1
XANTENNA__14677__A net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17500_ clknet_leaf_31_wb_clk_i _03187_ _01483_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09151__A1 _05490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1280 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1291 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2907 sky130_fd_sc_hd__dlygate4sd3_1
X_14712_ net1306 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11924_ net1883 _07941_ net481 vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15692_ net1219 vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14027__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17293__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ clknet_leaf_138_wb_clk_i _03118_ _01414_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14643_ net1247 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__inv_2
X_11855_ net2146 net305 net490 vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__mux2_1
X_18081__1581 vssd1 vssd1 vccd1 vccd1 _18081__1581/HI net1581 sky130_fd_sc_hd__conb_1
XFILLER_0_111_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10049__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17362_ clknet_leaf_129_wb_clk_i _03049_ _01345_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10806_ _07144_ _07145_ _07142_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14574_ net1337 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__inv_2
X_11786_ net1922 net309 net496 vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__mux2_1
XANTENNA__09454__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16313_ clknet_leaf_57_wb_clk_i _02067_ _00296_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13525_ net980 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _03979_ _03980_
+ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__a22o_1
XANTENNA__09002__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10737_ _06966_ _06967_ _06964_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__a21oi_1
X_17293_ clknet_leaf_2_wb_clk_i _02980_ _01276_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15301__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16244_ clknet_leaf_81_wb_clk_i _02004_ _00232_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13456_ _03914_ _03916_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10668_ net546 net373 _07007_ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ net2766 net234 net421 vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__mux2_1
XANTENNA__12136__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16175_ clknet_leaf_107_wb_clk_i _01935_ _00163_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10599_ net551 _06562_ vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10445__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13387_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _05727_ vssd1 vssd1
+ vccd1 vccd1 _03848_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10221__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
XFILLER_0_49_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
X_15126_ net1198 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
X_12338_ net2471 net237 net427 vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10772__A1 _06598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11975__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15057_ net1291 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12269_ net2730 net245 net435 vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__mux2_1
X_14008_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[57\] _04258_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[105\]
+ _04298_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_133_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09672__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11721__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09390__A1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__A _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15959_ net1406 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__inv_2
XANTENNA__10288__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ net730 _04752_ _04838_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09480_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[30\] net694 net663 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__a22o_1
XANTENNA__08585__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08431_ net1010 net920 vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__and2_2
X_17629_ clknet_leaf_111_wb_clk_i _03314_ _01570_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16660__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08362_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[30\] net743 _04681_
+ _04677_ _04670_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08293_ net1148 net1151 net1153 net1146 vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_117_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13529__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10460__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08751__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12046__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout303_A _07912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1045_A team_01_WB.instance_to_wrap.cpu.SR1.enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10212__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11885__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16040__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout301 _07921_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout312 net313 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09905__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout334 net335 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout672_A _04797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout345 _04748_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_2
XANTENNA__10802__B net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__B net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09381__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout356 _03741_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__dlymetal6s2s_1
X_09816_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\] net767 vssd1 vssd1
+ vccd1 vccd1 _06156_ sky130_fd_sc_hd__or2_1
Xfanout367 net368 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_2
Xfanout378 _04750_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__buf_4
Xfanout389 net390 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_8
XANTENNA__16190__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10521__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[20\] net745 _06072_
+ _06075_ _06076_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout937_A _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09678_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[22\] net815 net778 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__a22o_1
XANTENNA__14009__A2 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08629_ net600 _04968_ _04949_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11640_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _07817_ vssd1 vssd1
+ vccd1 vccd1 _07850_ sky130_fd_sc_hd__xor2_1
XANTENNA__09436__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11571_ net2700 net152 team_01_WB.instance_to_wrap.cpu.K0.next_state vssd1 vssd1
+ vccd1 vccd1 _03271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_64_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15121__A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13310_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] _07707_ vssd1 vssd1 vccd1 vccd1
+ _03792_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10522_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[31\] net889
+ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14290_ net1382 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10453_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[26\] net952
+ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__and3_1
X_13241_ net2784 net355 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1
+ vccd1 vccd1 _01909_ sky130_fd_sc_hd__a22o_1
XANTENNA__10265__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17509__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12743__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13172_ net134 net849 net841 net1751 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__a22o_1
X_10384_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[16\] net817 net779 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__a22o_1
XANTENNA_input66_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11795__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ net2355 net293 net456 vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__mux2_1
X_17980_ net1480 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_62_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12054_ net2254 net306 net466 vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__mux2_1
X_16931_ clknet_leaf_19_wb_clk_i _02618_ _00914_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16533__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ _05729_ _06812_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__and2_1
X_16862_ clknet_leaf_44_wb_clk_i _02549_ _00845_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15813_ net1310 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__inv_2
Xfanout890 net891 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__buf_4
XFILLER_0_137_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16793_ clknet_leaf_46_wb_clk_i _02480_ _00776_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11824__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15744_ net1238 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12956_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[4\] _05110_ net1034 vssd1
+ vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__mux2_2
XFILLER_0_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11907_ net1810 net267 net479 vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13208__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15675_ net1183 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__inv_2
X_12887_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[26\] _03665_ net1030 vssd1
+ vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17414_ clknet_leaf_41_wb_clk_i _03101_ _01397_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14626_ net1205 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17039__CLK clknet_leaf_143_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11838_ net2906 net271 net488 vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09427__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17345_ clknet_leaf_48_wb_clk_i _03032_ _01328_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14557_ net1406 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11769_ net2928 net243 net495 vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13508_ net726 _07056_ net981 vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__a21oi_1
X_17276_ clknet_leaf_37_wb_clk_i _02963_ _01259_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14488_ net1330 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__inv_2
XANTENNA__09667__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10993__A1 _05115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_0__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__08571__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16227_ clknet_leaf_105_wb_clk_i net1944 _00215_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
XANTENNA__16063__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17189__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13439_ _03883_ _03896_ _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12734__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16158_ clknet_leaf_101_wb_clk_i _01921_ _00146_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15109_ net1209 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__inv_2
X_08980_ _05307_ _05311_ _05315_ _05319_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__and4bb_1
X_16089_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[11\]
+ _00077_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10840__S1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08299__B net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10341__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09601_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[24\] net952
+ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09532_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[28\] net973
+ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08746__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] net713 _04841_ vssd1 vssd1
+ vccd1 vccd1 _05803_ sky130_fd_sc_hd__a21o_1
XANTENNA__08874__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout253_A _07904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08414_ net712 _04751_ _04752_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__nor3_4
XANTENNA__10681__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09394_ net560 _05659_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08345_ net988 net954 vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__and2_1
XANTENNA__12422__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08626__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16406__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout420_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1162_A team_01_WB.instance_to_wrap.cpu.f0.state\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08276_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] net2047 net1037 vssd1 vssd1
+ vccd1 vccd1 _03411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16556__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13396__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout887_A _04799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12504__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18080__1580 vssd1 vssd1 vccd1 vccd1 _18080__1580/HI net1580 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_110_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1107 net1108 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__buf_1
XFILLER_0_121_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1118 net1127 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__buf_2
Xfanout1129 net1135 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_111_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout186 _07639_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_2
XFILLER_0_138_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_2
XANTENNA__13843__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12810_ net1728 net641 net608 _03635_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__a22o_1
X_13790_ net1170 _04160_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[28\] _07088_ net1026 vssd1 vssd1
+ vccd1 vccd1 _03588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15460_ net1237 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__inv_2
X_12672_ net2729 net261 net388 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14411_ net1360 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__inv_2
X_11623_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[27\] _07566_ net715 vssd1 vssd1
+ vccd1 vccd1 _07836_ sky130_fd_sc_hd__mux2_1
XANTENNA__08617__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15391_ net1254 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17331__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17130_ clknet_leaf_11_wb_clk_i _02817_ _01113_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14342_ net1373 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11554_ net37 net36 net35 net34 vssd1 vssd1 vccd1 vccd1 _07786_ sky130_fd_sc_hd__nor4_1
XFILLER_0_110_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17061_ clknet_leaf_31_wb_clk_i _02748_ _01044_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10505_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[31\] net760 net755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__a22o_1
X_14273_ net1368 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[20\] net579 vssd1 vssd1 vccd1
+ vccd1 _07770_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16012_ net1385 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13224_ net2672 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1
+ vccd1 vccd1 _01926_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10436_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[27\] net741 _06774_ _06775_
+ net770 vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__a2111o_1
X_13155_ net1943 net843 net840 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[21\] vssd1
+ vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a22o_1
XANTENNA__12414__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10367_ net581 _06706_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] net626
+ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__a2bb2o_4
X_12106_ net1850 net267 net456 vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__mux2_1
X_17963_ net1463 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_104_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13086_ net2410 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[8\] net860 vssd1 vssd1
+ vccd1 vccd1 _02039_ sky130_fd_sc_hd__mux2_1
X_10298_ net559 _04919_ _05731_ _06637_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_40_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13141__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16914_ clknet_leaf_132_wb_clk_i _02601_ _00897_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12037_ net2505 net272 net465 vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__mux2_1
X_17894_ net1597 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XANTENNA__09896__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16845_ clknet_leaf_140_wb_clk_i _02532_ _00828_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16776_ clknet_leaf_21_wb_clk_i _02463_ _00759_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13988_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[88\] _04241_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[120\]
+ _04270_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09648__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08566__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15727_ net1217 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__inv_2
XANTENNA__08856__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ net2488 net871 net358 _03702_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16429__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15658_ net1282 vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08863__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14609_ net1365 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15589_ net1210 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08130_ team_01_WB.instance_to_wrap.cpu.f0.i\[30\] _04493_ team_01_WB.instance_to_wrap.cpu.f0.num\[7\]
+ _04486_ _04582_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17328_ clknet_leaf_15_wb_clk_i _03015_ _01311_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12955__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16579__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14157__A1 _04195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08061_ _04522_ _04528_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_133_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17259_ clknet_leaf_2_wb_clk_i _02946_ _01242_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09694__A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10194__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08963_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] net595 vssd1 vssd1 vccd1
+ vccd1 _05303_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13132__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08894_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[2\] net928 vssd1
+ vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__and3_1
XANTENNA__10071__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1008_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17204__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout370_A net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14093__B1 _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08476__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09515_ _05851_ _05852_ _05853_ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14775__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17354__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1377_A net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10654__A0 _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09446_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[29\] net916 vssd1
+ vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08773__A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13199__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout802_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[26\] net663 net650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[26\]
+ _05714_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12946__A2 _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08328_ net1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[30\] net969
+ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10957__A1 _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09811__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1652_A team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09100__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ net1779 net2562 net1037 vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11270_ _07605_ _07608_ _07609_ vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10709__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10221_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] net767 net623 vssd1
+ vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12234__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10543__A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[11\] net744 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[11\]
+ _06491_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__a221o_1
XANTENNA__13659__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13123__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14960_ net1272 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__inv_2
X_10083_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[7\] net772 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[7\]
+ _06416_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__a221o_1
XANTENNA__08948__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[22\] vssd1 vssd1 vccd1 vccd1 net1625
+ sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\] _04207_ vssd1 vssd1 vccd1
+ vccd1 _04209_ sky130_fd_sc_hd__and2_1
X_14891_ net1296 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16630_ clknet_leaf_0_wb_clk_i _02317_ _00613_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13842_ net1165 net1061 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[3\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[3\] sky130_fd_sc_hd__and3b_1
XANTENNA__10893__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14084__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16561_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[27\]
+ _00544_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13773_ _04154_ _04158_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11437__A2 _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ net547 _06398_ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_84_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10645__A0 _06098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15512_ net1179 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12724_ net1027 _03573_ _03574_ net1161 vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__a211o_1
X_16492_ clknet_leaf_108_wb_clk_i _02246_ _00475_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15443_ net1278 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12655_ net2959 net189 net389 vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12409__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11606_ _07796_ _07822_ net614 vssd1 vssd1 vccd1 vccd1 _07823_ sky130_fd_sc_hd__mux2_2
XANTENNA__13595__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15374_ net1283 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_122_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12586_ net1896 net314 net401 vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__mux2_1
XANTENNA__09263__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09802__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17113_ clknet_leaf_55_wb_clk_i _02800_ _01096_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14325_ net1356 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__inv_2
X_18093_ net1587 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
X_11537_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[16\] net1157 net587 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__a22o_1
XANTENNA__09010__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold409 team_01_WB.instance_to_wrap.a1.ADR_I\[22\] vssd1 vssd1 vccd1 vccd1 net2025
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17044_ clknet_leaf_13_wb_clk_i _02731_ _01027_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output97_A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14256_ net1323 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__inv_2
X_11468_ net368 _07761_ net3001 net875 vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_81_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13207_ net32 net837 net630 net2424 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__a22o_1
X_10419_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[27\] net952
+ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__and3b_1
X_14187_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\]
+ _04453_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12144__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10176__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ team_01_WB.instance_to_wrap.cpu.f0.i\[25\] _07695_ vssd1 vssd1 vccd1 vccd1
+ _07723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13138_ net102 net850 net633 net1650 vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__a22o_1
XANTENNA__11983__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13069_ net2875 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[25\] net866 vssd1 vssd1
+ vccd1 vccd1 _02056_ sky130_fd_sc_hd__mux2_1
X_17946_ net1446 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
Xhold1109 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[106\] vssd1 vssd1 vccd1 vccd1
+ net2725 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_131_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08858__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09869__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17877_ clknet_leaf_99_wb_clk_i net1642 _01817_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11284__A _07135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16828_ clknet_leaf_36_wb_clk_i _02515_ _00811_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14075__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11428__A2 _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16759_ clknet_leaf_138_wb_clk_i _02446_ _00742_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09300_ net1073 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[22\] net878
+ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__and3_1
XANTENNA__10636__A0 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09231_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[21\] net886 vssd1
+ vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_1499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12319__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12928__A2 _07757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09162_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[16\] net928
+ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__and3_1
XANTENNA__08057__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08113_ team_01_WB.instance_to_wrap.cpu.f0.i\[29\] team_01_WB.instance_to_wrap.cpu.f0.num\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09093_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[13\] net920 vssd1
+ vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout216_A _07835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08044_ net1927 net570 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1
+ vccd1 vccd1 _03547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold910 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold921 _03525_ vssd1 vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold932 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[22\] vssd1 vssd1 vccd1 vccd1 net2548
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09557__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold943 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold954 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12054__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10167__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1125_A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold965 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[102\] vssd1 vssd1 vccd1 vccd1
+ net2592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 team_01_WB.instance_to_wrap.cpu.f0.num\[11\] vssd1 vssd1 vccd1 vccd1 net2603
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09995_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[2\] net776 net738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__a22o_1
XANTENNA__12989__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout585_A net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[6\] net890 vssd1
+ vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_4_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1610 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1621 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1632 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3248 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[3\] net676 net661 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[3\]
+ net707 vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1643 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3259 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10810__B _05261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout752_A _04678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1654 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 net3270
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08532__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1665 team_01_WB.instance_to_wrap.a1.ADR_I\[10\] vssd1 vssd1 vccd1 vccd1 net3281
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1676 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 net3292
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10088__D1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09599__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ _07103_ _07109_ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08934__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09429_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[28\] net668 net667 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[28\]
+ _05768_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_118_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12229__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16894__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12440_ net2388 net233 net416 vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08599__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12371_ net1842 net236 net423 vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__mux2_1
XANTENNA__13592__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14110_ _04217_ _04231_ _04239_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__and3_1
X_11322_ _07657_ net1960 _07655_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__mux2_1
XANTENNA__16124__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15090_ net1231 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14041_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[75\] _04268_ _04289_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__a22o_1
X_11253_ _07055_ _07278_ vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10273__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10158__A2 _05379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10204_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[8\] net941 vssd1
+ vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__and3_1
X_11184_ _07014_ _07149_ _07242_ net525 vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__a22o_1
X_17800_ clknet_leaf_65_wb_clk_i net2513 _01740_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[70\]
+ sky130_fd_sc_hd__dfrtp_1
X_10135_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[11\] net793 net753 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[11\]
+ _06473_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15992_ net1336 vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13501__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ _06404_ _06405_ _06316_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__a21oi_2
X_17731_ clknet_leaf_81_wb_clk_i _03407_ _01671_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14943_ net1255 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__inv_2
XANTENNA__11658__A2 _07171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17662_ clknet_leaf_114_wb_clk_i _03347_ _01603_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14874_ net1186 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
XANTENNA__10330__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16613_ clknet_leaf_31_wb_clk_i _02300_ _00596_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_82_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13825_ net2459 net831 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[18\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_67_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17593_ clknet_leaf_69_wb_clk_i _03280_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09005__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16544_ clknet_leaf_112_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[10\]
+ _00527_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13756_ _04143_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__nor2_1
X_10968_ _07276_ _07306_ _07307_ _07299_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__o211a_2
X_12707_ net2550 net289 net385 vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__mux2_1
XANTENNA__11551__B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09302__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16475_ clknet_leaf_84_wb_clk_i _02229_ _00458_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11291__B1 _06960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10448__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13687_ team_01_WB.instance_to_wrap.cpu.c0.count\[15\] _04109_ vssd1 vssd1 vccd1
+ vccd1 _04110_ sky130_fd_sc_hd__or2_1
XANTENNA__12139__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10899_ net555 _07238_ _06963_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_14_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13568__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15426_ net1264 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12638_ net2751 net232 net394 vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11978__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15357_ net1253 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__inv_2
XANTENNA__13583__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ net2580 net237 net399 vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10397__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14308_ net1350 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__inv_2
XANTENNA__12791__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18076_ net1576 vssd1 vssd1 vccd1 vccd1 la_data_out[118] sky130_fd_sc_hd__buf_2
X_15288_ net1171 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__inv_2
Xhold206 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 _02151_ vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09675__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold228 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
X_17027_ clknet_leaf_19_wb_clk_i _02714_ _01010_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold239 team_01_WB.instance_to_wrap.cpu.RU0.state\[2\] vssd1 vssd1 vccd1 vccd1 net1855
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ net1352 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10149__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout708 net709 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_2
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout719 _04723_ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_124_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[0\] net663 _05138_ _05139_
+ net709 vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_52_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08762__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12602__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[15\] net758 net737 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[5\] net690 _05057_ _05058_
+ _05063_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__a2111o_1
X_17929_ net1431 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_20_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10630__B net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1290 net1294 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__buf_2
XANTENNA__10857__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08662_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[10\] net696 _04973_
+ _04976_ net706 vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__a2111o_1
XANTENNA_clkbuf_leaf_89_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14048__B1 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08593_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[15\] net654 _04921_
+ _04924_ _04927_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10609__A0 _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08754__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09212__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12049__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1075_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13559__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[17\] _04776_ _05541_
+ _05546_ _05551_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11888__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09145_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[14\] net674 _05470_ _05474_
+ _05478_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13574__A2 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout500_A _07795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1242_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10388__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09242__A3 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09076_ _05380_ _05415_ net602 vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__mux2_2
XFILLER_0_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08027_ _04512_ _04522_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__nor2_4
Xhold740 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11337__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold751 team_01_WB.instance_to_wrap.cpu.f0.num\[16\] vssd1 vssd1 vccd1 vccd1 net2367
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09882__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold784 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 _02039_ vssd1 vssd1 vccd1 vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_89_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12512__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ net993 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[2\] net955 vssd1
+ vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_18_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08929__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[6\] net887 vssd1
+ vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__and3_1
XANTENNA__17692__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1440 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1451 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11940_ net2172 net268 net475 vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14039__B1 _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1462 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1473 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10312__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1484 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[24\] vssd1 vssd1 vccd1 vccd1
+ net3100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1495 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3111 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13851__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11871_ net1932 net273 net485 vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13610_ _03883_ _03895_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08269__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10822_ net553 _07160_ _07161_ _06964_ vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14590_ net1337 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09122__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13541_ net197 net193 _07854_ net643 vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__o211a_1
XANTENNA__11371__B team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10753_ _06034_ _07091_ _06001_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14963__A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16260_ clknet_leaf_104_wb_clk_i net2026 _00248_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
X_13472_ _03924_ _03929_ _03932_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17072__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ net540 _07022_ _06970_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_47_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ net1298 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11798__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ _07942_ _07946_ net573 vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__and3_4
X_16191_ clknet_leaf_115_wb_clk_i _01951_ _00179_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13565__A2 _07135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10379__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15142_ net1324 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12354_ net3014 net320 net430 vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__mux2_1
XANTENNA__13298__B net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10715__B _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11305_ net727 _07476_ net187 _07644_ vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__a22o_1
XANTENNA__13317__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15073_ net1200 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__inv_2
X_12285_ net1964 net294 net438 vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14024_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[74\] _04235_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09792__A _06129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11236_ _06906_ _07027_ _07033_ _05263_ net339 vssd1 vssd1 vccd1 vccd1 _07576_ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_123_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11167_ _07502_ _07506_ _07494_ vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__and3b_2
XFILLER_0_101_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10731__A _05115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12422__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10118_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[6\] net814 _04659_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[6\]
+ _06444_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_69_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ net1409 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__inv_2
X_11098_ _07431_ _07437_ _07339_ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_69_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17714_ clknet_leaf_81_wb_clk_i _03398_ _01655_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14926_ net1284 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
X_10049_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[0\] net775 net746 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10303__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17645_ clknet_leaf_111_wb_clk_i _03330_ _01586_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\]
+ sky130_fd_sc_hd__dfrtp_4
X_14857_ net1215 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_118_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13808_ net2066 net833 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[1\]
+ sky130_fd_sc_hd__and2_1
X_17576_ clknet_leaf_72_wb_clk_i _03263_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dfxtp_1
X_14788_ net1306 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__inv_2
XANTENNA__09457__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08574__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16527_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[25\]
+ _00510_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13739_ net3004 _04524_ team_01_WB.instance_to_wrap.cpu.f0.next_lcd_en vssd1 vssd1
+ vccd1 vccd1 _00024_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16458_ clknet_leaf_139_wb_clk_i _02212_ _00441_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15409_ net1288 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__inv_2
X_16389_ clknet_leaf_76_wb_clk_i net2535 _00372_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10625__B net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18059_ net1559 vssd1 vssd1 vccd1 vccd1 la_data_out[101] sky130_fd_sc_hd__buf_2
XFILLER_0_44_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09901_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[5\] net780 net742 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__a22o_1
XANTENNA__10344__C net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout505 _06636_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__buf_2
Xfanout516 _05261_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09832_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[13\] net807 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[13\]
+ _06171_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__a221o_1
Xfanout527 _05223_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_2
Xfanout538 net539 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12332__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout549 _05151_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08749__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09207__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ _06000_ _06034_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__nand2_1
XANTENNA__08111__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[5\] net883 vssd1
+ vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09694_ net509 _06033_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__and2_1
X_17959__1459 vssd1 vssd1 vccd1 vccd1 _17959__1459/HI net1459 sky130_fd_sc_hd__conb_1
XFILLER_0_136_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08645_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[10\] net909
+ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout450_A _07958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1192_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08576_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[19\] net698 _04913_
+ _04914_ _04915_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09448__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13244__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17095__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10058__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08484__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09999__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_136_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_136_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout715_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire917 net918 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13399__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12507__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09128_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[14\] net888
+ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__and3_1
XANTENNA__09620__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16932__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09059_ net1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[12\] net880
+ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12070_ net2683 net271 net461 vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__mux2_1
XANTENNA__13846__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold570 team_01_WB.instance_to_wrap.cpu.f0.num\[4\] vssd1 vssd1 vccd1 vccd1 net2186
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12750__B net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold592 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08726__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11021_ _07360_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__inv_2
XANTENNA__12242__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10533__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11366__B team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15760_ net1401 vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__inv_2
X_12972_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[114\] net1904 net868 vssd1 vssd1
+ vccd1 vccd1 _02153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09687__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1270 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[25\] vssd1 vssd1 vccd1 vccd1
+ net2886 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ net2916 net314 net482 vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14711_ net1304 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__inv_2
Xhold1281 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2897 sky130_fd_sc_hd__dlygate4sd3_1
X_15691_ net1298 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__inv_2
XANTENNA__11494__B1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1292 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14642_ net1223 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ clknet_leaf_1_wb_clk_i _03117_ _01413_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11854_ net3130 net310 net489 vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13235__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_95_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10805_ _05657_ net332 _07143_ net337 net370 vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__a221o_1
X_14573_ net1409 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17361_ clknet_leaf_14_wb_clk_i _03048_ _01344_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11785_ net1965 net297 net497 vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16312_ clknet_leaf_73_wb_clk_i _02066_ _00295_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_13524_ net722 _07588_ net1066 vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17292_ clknet_leaf_130_wb_clk_i _02979_ _01275_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10736_ _07074_ _07075_ _07072_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_138_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16243_ clknet_leaf_81_wb_clk_i net1651 _00231_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13455_ _03859_ _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__and2b_1
XFILLER_0_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10667_ net552 _06250_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__nor2_1
XANTENNA__12417__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12746__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12406_ net2666 net264 net420 vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13102__A net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16174_ clknet_leaf_107_wb_clk_i _01934_ _00162_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09072__D1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13386_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _05757_ vssd1 vssd1
+ vccd1 vccd1 _03847_ sky130_fd_sc_hd__and2_1
XANTENNA__09611__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10598_ _06936_ _06937_ net539 vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__mux2_1
XANTENNA__10221__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15125_ net1221 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__inv_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
X_12337_ net2076 net239 net427 vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__mux2_1
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12941__A team_01_WB.instance_to_wrap.cpu.f0.write_data\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10164__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10772__A2 _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15056_ net1226 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__inv_2
X_12268_ net2644 net203 net435 vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__mux2_1
XANTENNA__13171__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14007_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[33\] _04230_ _04240_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[89\]
+ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11219_ _05758_ _07558_ vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__nand2_1
XANTENNA__12152__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11958__A_N team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12199_ net2407 net205 net443 vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__mux2_1
XANTENNA__11182__C1 _06915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10524__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XANTENNA__08569__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09390__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11991__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15958_ net1392 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13474__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09678__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08866__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13474__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09142__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14909_ net1250 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15889_ net1337 vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08350__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08430_ net1109 net1112 net1114 net1106 vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__and4bb_2
X_17628_ clknet_leaf_110_wb_clk_i _03313_ _01569_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13226__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15699__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08361_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[30\] net819 net807 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17559_ clknet_leaf_138_wb_clk_i _03246_ _01542_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10339__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08292_ net1128 net975 vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__and2_2
XFILLER_0_116_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09850__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12327__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12737__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1038_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10074__C net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13162__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_2
XFILLER_0_100_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout313 _07931_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12062__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1205_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout335 _06918_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout346 net348 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_4
X_09815_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[14\] net817 net762 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[14\]
+ _06154_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__a221o_1
Xfanout357 net358 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_2
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12997__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout368 _07759_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_2
Xfanout379 net382 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_8
XANTENNA_fanout665_A _04806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[20\] net813 _06074_ _06079_
+ _06082_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__a2111o_1
X_09677_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[22\] net756 _06005_ _06007_
+ _06015_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout832_A team_01_WB.instance_to_wrap.cpu.RU0.next_ihit vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08628_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\] net705 _04961_ _04967_
+ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__o22a_4
XFILLER_0_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09728__A_N net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08559_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[19\] net685 _04896_
+ _04897_ _04898_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_33_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10436__D1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11570_ team_01_WB.instance_to_wrap.cpu.K0.count\[1\] team_01_WB.instance_to_wrap.cpu.K0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__or2_1
XFILLER_0_33_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09841__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08942__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10521_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[31\] net934 vssd1
+ vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__and3_1
XANTENNA__17880__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12237__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13240_ net2202 net356 net352 team_01_WB.instance_to_wrap.cpu.f0.i\[10\] vssd1 vssd1
+ vccd1 vccd1 _01910_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10452_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[26\] net964
+ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13171_ net135 net849 net841 net1837 vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10383_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[16\] net798 net788 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[16\]
+ _06722_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17110__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12122_ net2873 net316 net458 vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_33_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input59_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13153__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11377__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16930_ clknet_leaf_35_wb_clk_i _02617_ _00913_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12053_ net1901 net309 net463 vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18109__1592 vssd1 vssd1 vccd1 vccd1 _18109__1592/HI net1592 sky130_fd_sc_hd__conb_1
XANTENNA__10506__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11703__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ _07342_ _07343_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__or2_1
XANTENNA__09372__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16861_ clknet_leaf_49_wb_clk_i _02548_ _00844_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout880 _04810_ vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__buf_4
XANTENNA__08580__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15812_ net1310 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__inv_2
Xfanout891 _04796_ vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__buf_4
XANTENNA__12700__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16792_ clknet_leaf_27_wb_clk_i _02479_ _00775_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12955_ net1837 net872 net359 _03712_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a22o_1
X_15743_ net1256 vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__inv_2
XANTENNA__11824__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11906_ net1785 net236 net479 vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__mux2_1
X_18029__1529 vssd1 vssd1 vccd1 vccd1 _18029__1529/HI net1529 sky130_fd_sc_hd__conb_1
XANTENNA__08883__A1 _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15674_ net1190 vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__inv_2
X_12886_ _05726_ net577 net361 vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__o21ba_1
XANTENNA__16978__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17413_ clknet_leaf_39_wb_clk_i _03100_ _01396_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14625_ net1366 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__inv_2
X_11837_ net3157 net244 net487 vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__mux2_1
XANTENNA__09013__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14556_ net1392 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__inv_2
X_17344_ clknet_leaf_33_wb_clk_i _03031_ _01327_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11768_ net3194 net201 net495 vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__mux2_1
XANTENNA__09832__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09948__C _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08852__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16208__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10719_ _07001_ _07008_ net534 vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__mux2_1
X_13507_ net186 _03964_ _03965_ net726 vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14487_ net1332 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__inv_2
XANTENNA__12147__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17275_ clknet_leaf_50_wb_clk_i _02962_ _01258_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11699_ net1958 net289 net502 vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16226_ clknet_leaf_104_wb_clk_i net2309 _00214_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13438_ _03889_ _03891_ _03897_ _03898_ _03885_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__o32a_1
XANTENNA__12195__A1 _07838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11986__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16157_ clknet_leaf_97_wb_clk_i _01920_ _00145_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_17958__1458 vssd1 vssd1 vccd1 vccd1 _17958__1458/HI net1458 sky130_fd_sc_hd__conb_1
XFILLER_0_49_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13369_ net585 net564 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1
+ vccd1 _03837_ sky130_fd_sc_hd__o21a_1
XANTENNA__16358__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15108_ net1193 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__inv_2
X_16088_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[10\]
+ _00076_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11287__A _06961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15982__A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15039_ net1254 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09600_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[24\] net806 net777 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__a22o_1
XANTENNA__12610__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09531_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[28\] net969
+ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09462_ _05788_ _05791_ _05801_ net704 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__o32a_2
XFILLER_0_66_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08413_ net720 _04751_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09393_ _05570_ _05620_ _05658_ net559 vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout246_A _07862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08344_ net990 net943 vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__and2_4
XFILLER_0_30_1626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08275_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[6\] net1960 net1037 vssd1 vssd1
+ vccd1 vccd1 _03412_ sky130_fd_sc_hd__mux2_1
XANTENNA__12057__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17133__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout413_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13099__D _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11896__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1322_A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17283__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout782_A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13135__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1108 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[23\] vssd1 vssd1 vccd1 vccd1
+ net1108 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1119 net1127 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09890__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09354__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout187 net188 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12520__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout198 _07633_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09106__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09729_ _06066_ _06067_ net508 vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__a21boi_1
XANTENNA__11449__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13989__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12740_ net1790 net639 net606 _03587_ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12671_ net2820 net231 net389 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14410_ net1338 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__inv_2
XANTENNA__15132__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11622_ net3120 net216 net499 vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__mux2_1
X_15390_ net1251 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__inv_2
XANTENNA__09814__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08672__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09130__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14341_ net1370 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__inv_2
X_11553_ net2491 net1160 net589 vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10975__A2 _06465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17060_ clknet_leaf_51_wb_clk_i _02747_ _01043_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10504_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[31\] net808 net758 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[31\]
+ _06832_ vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14272_ net1367 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__inv_2
X_11484_ net367 _07769_ net1918 net875 vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_68_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16500__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16011_ net1385 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__inv_2
X_13223_ net3074 net353 net349 net1062 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10435_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[27\] net803 _06752_
+ _06753_ _06754_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11924__A1 _07941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13154_ net1707 net843 net840 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[22\] vssd1
+ vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10366_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] net765 net622 vssd1
+ vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13126__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12105_ net2845 net236 net455 vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__mux2_1
X_17962_ net1462 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
X_13085_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\] net2727 net868 vssd1 vssd1
+ vccd1 vccd1 _02040_ sky130_fd_sc_hd__mux2_1
XANTENNA__16650__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10297_ _04883_ _05568_ _04919_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_97_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12036_ net3229 net245 net464 vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__mux2_1
X_16913_ clknet_leaf_15_wb_clk_i _02600_ _00896_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_17893_ net1596 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XANTENNA__09008__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16844_ clknet_leaf_133_wb_clk_i _02531_ _00827_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12430__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14211__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10360__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16775_ clknet_leaf_16_wb_clk_i _02462_ _00758_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13987_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[64\] _04233_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[120\]
+ _04278_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15726_ net1284 vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__inv_2
XANTENNA__10112__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12938_ _03694_ _03701_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[11\] net1028
+ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15657_ net1229 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__inv_2
X_12869_ _06881_ net577 net361 vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_56_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15042__A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14608_ net1330 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__inv_2
XANTENNA__13601__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09805__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15588_ net1238 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08582__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17327_ clknet_leaf_144_wb_clk_i _03014_ _01310_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14539_ net1408 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10966__A2 _06921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08060_ _04522_ _04532_ _04536_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__o21bai_1
XANTENNA_wire583_A _05040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17258_ clknet_leaf_3_wb_clk_i _02945_ _01241_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16209_ clknet_leaf_78_wb_clk_i net1694 _00197_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10179__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17189_ clknet_leaf_31_wb_clk_i _02876_ _01172_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12605__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09584__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13117__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08962_ _05043_ _05301_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09336__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08893_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[2\] net939 vssd1
+ vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_127_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11745__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12340__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10351__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12891__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14093__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09514_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[29\] net801 net786 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[29\] net939
+ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10654__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout530_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08773__B _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09376_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[26\] net688 net673 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[26\]
+ _05715_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_1600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10406__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08327_ net1134 net969 vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__and2_4
XANTENNA__15887__A net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09885__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14148__A2 _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08258_ net3015 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[15\] net1047 vssd1 vssd1
+ vccd1 vccd1 _03429_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout997_A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12515__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16673__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08189_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[92\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[84\]
+ net1041 vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10220_ _06550_ _06552_ _06556_ _06559_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__or4_4
XFILLER_0_42_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09575__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13108__A0 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10543__B _06882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18028__1528 vssd1 vssd1 vccd1 vccd1 _18028__1528/HI net1528 sky130_fd_sc_hd__conb_1
XFILLER_0_24_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10151_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[11\] net790 net742 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17029__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09327__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13854__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[7\] net739 _06412_ _06418_
+ _06419_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__a2111o_1
X_13910_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\] _04207_ vssd1 vssd1 vccd1
+ vccd1 _04208_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12250__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14890_ net1279 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08667__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ net1165 net1061 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[2\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[2\] sky130_fd_sc_hd__and3b_1
XFILLER_0_138_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17179__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13772_ _04156_ _01836_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__or2_1
X_16560_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[26\]
+ _00543_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10984_ _07277_ _07283_ net526 vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__mux2_1
XANTENNA__08964__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957__1457 vssd1 vssd1 vccd1 vccd1 _17957__1457/HI net1457 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_84_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10645__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15511_ net1196 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__inv_2
X_12723_ net1027 team_01_WB.instance_to_wrap.cpu.f0.write_i vssd1 vssd1 vccd1 vccd1
+ _03574_ sky130_fd_sc_hd__nor2_1
X_16491_ clknet_leaf_104_wb_clk_i _02245_ _00474_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15442_ net1232 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12654_ _07791_ _07793_ net573 vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11605_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] _07821_ vssd1 vssd1
+ vccd1 vccd1 _07822_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_61_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ net3265 net319 net402 vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__mux2_1
X_15373_ net1213 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17112_ clknet_leaf_30_wb_clk_i _02799_ _01095_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14139__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11536_ net2170 net1157 net587 net1150 vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__a22o_1
X_14324_ net1356 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__inv_2
XANTENNA__11070__B2 _04969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18092_ net637 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13347__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17043_ clknet_leaf_135_wb_clk_i _02730_ _01026_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14255_ net1323 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_78_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11467_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[29\] net580 vssd1 vssd1 vccd1
+ vccd1 _07761_ sky130_fd_sc_hd__nand2_1
XANTENNA__12425__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10734__A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13206_ net33 net836 net629 net1672 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__o22a_1
X_10418_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[27\] net944
+ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__and3b_1
X_14186_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\] _04453_ net1987 vssd1
+ vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11549__B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11398_ _04468_ _07721_ _07722_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13137_ net103 net850 net633 net3125 vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10349_ net987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[17\] net966 vssd1
+ vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__and3_1
X_13068_ net2566 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[26\] net858 vssd1 vssd1
+ vccd1 vccd1 _02057_ sky130_fd_sc_hd__mux2_1
X_17945_ net1445 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XANTENNA__12322__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ net1928 net295 net468 vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__mux2_1
XANTENNA__12160__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_79_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17876_ clknet_leaf_97_wb_clk_i _03551_ _01816_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16827_ clknet_leaf_17_wb_clk_i _02514_ _00810_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11284__B _07611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10884__A1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10884__B2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16758_ clknet_leaf_140_wb_clk_i _02445_ _00741_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10636__A1 _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15709_ net1251 vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__inv_2
X_16689_ clknet_leaf_18_wb_clk_i _02376_ _00672_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_09230_ net377 net343 _05493_ _05569_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__and4_2
XANTENNA__11079__A_N net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12389__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09161_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[16\] net924
+ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08057__A2 team_01_WB.instance_to_wrap.cpu.K0.keyvalid vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09254__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09201__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08112_ _04480_ team_01_WB.instance_to_wrap.cpu.f0.num\[14\] team_01_WB.instance_to_wrap.cpu.f0.num\[9\]
+ _04484_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a22o_1
XANTENNA__10347__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09092_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[13\] net881 vssd1
+ vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08043_ net2398 net570 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1
+ vccd1 vccd1 _03548_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12335__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold900 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold911 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout209_A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold933 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[40\] vssd1 vssd1 vccd1 vccd1
+ net2560 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08114__A team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold955 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09994_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[2\] net816 net813 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1020_A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1118_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09309__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08945_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[6\] net898 vssd1
+ vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout480_A _07949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1600 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3216 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12070__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1611 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3227 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08876_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[3\] _04771_ _05199_ _05203_
+ _05205_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_4_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1622 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[23\] vssd1 vssd1 vccd1 vccd1
+ net3238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1633 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1644 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09319__A_N _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3271 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09190__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1666 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 net3282
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14786__A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout745_A _04684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout912_A _04779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10819__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09428_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[28\] net663 net649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09359_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[25\] net690 net687 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__a22o_1
XANTENNA__08048__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15410__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09796__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12370_ net1813 net241 net423 vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13849__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13329__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11321_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\] net1162 _04534_ _07652_ vssd1
+ vssd1 vccd1 vccd1 _07657_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12245__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14040_ net147 net604 vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11252_ _05681_ _06919_ net511 vssd1 vssd1 vccd1 vccd1 _07592_ sky130_fd_sc_hd__or3b_1
XFILLER_0_120_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11369__B _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[8\] net947 vssd1
+ vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_73_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_113_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11183_ net338 _07376_ _07522_ vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10134_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[11\] net967
+ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__and3_1
XANTENNA_input41_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15991_ net1405 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17730_ clknet_leaf_82_wb_clk_i _03406_ _01670_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10065_ _06313_ _06315_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__xor2_1
X_14942_ net1275 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__inv_2
XANTENNA__10866__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09720__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17661_ clknet_leaf_120_wb_clk_i _03346_ _01602_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10866__B2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14873_ net1258 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16612_ clknet_leaf_53_wb_clk_i _02299_ _00595_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13824_ net2080 net831 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[17\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_67_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17592_ clknet_leaf_69_wb_clk_i _03279_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13265__C1 _04466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16543_ clknet_leaf_112_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[9\]
+ _00526_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13755_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__or4b_1
X_10967_ net344 _07294_ _07305_ _07071_ vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__o22a_1
XANTENNA__10729__A _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12706_ net2318 net255 net384 vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10094__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16474_ clknet_leaf_82_wb_clk_i _02228_ _00457_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10898_ net528 _07237_ _07235_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__a21boi_1
X_13686_ team_01_WB.instance_to_wrap.cpu.c0.count\[14\] team_01_WB.instance_to_wrap.cpu.c0.count\[13\]
+ _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_14_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15425_ net1246 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__inv_2
XANTENNA__09021__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12637_ net2811 net264 net391 vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08039__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13742__A_N net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15356_ net1171 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__inv_2
X_12568_ net1864 net241 net399 vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__mux2_1
XANTENNA__09956__C net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08860__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12791__A1 team_01_WB.instance_to_wrap.a1.ADR_I\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_135_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14307_ net1357 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__inv_2
X_11519_ team_01_WB.instance_to_wrap.cpu.DM0.enable net717 vssd1 vssd1 vccd1 vccd1
+ _07783_ sky130_fd_sc_hd__nor2_1
XANTENNA__12155__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18075_ net1575 vssd1 vssd1 vccd1 vccd1 la_data_out[117] sky130_fd_sc_hd__buf_2
XFILLER_0_48_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15287_ net1196 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__inv_2
X_12499_ net2582 net201 net407 vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold207 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[3\] vssd1 vssd1 vccd1 vccd1
+ net1834 sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ clknet_leaf_33_wb_clk_i _02713_ _01009_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold229 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ net1367 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11994__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14169_ net1936 _04189_ _04445_ net1412 vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__a211oi_1
Xfanout709 _04757_ vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__buf_4
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[5\] net677 _05060_ net707
+ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_33_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11295__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17928_ net1616 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
XFILLER_0_59_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1280 net1286 vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__buf_4
X_08661_ _04997_ _04998_ _04999_ _05000_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__or4_1
XANTENNA__10857__A1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1291 net1293 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__buf_4
XANTENNA__09711__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17494__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10857__B2 _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17859_ clknet_leaf_90_wb_clk_i _03534_ _01799_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.read_i
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08592_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[15\] net686 _04808_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[15\] vssd1 vssd1 vccd1 vccd1
+ _04932_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10609__A1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10639__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18027__1527 vssd1 vssd1 vccd1 vccd1 _18027__1527/HI net1527 sky130_fd_sc_hd__conb_1
XFILLER_0_76_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10085__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08109__A _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09213_ net1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[17\] net882
+ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout326_A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10077__C net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[14\] net684 _05464_
+ _05466_ _05471_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_96_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1068_A team_01_WB.instance_to_wrap.cpu.IM0.pc_enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09075_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\] net705 _05411_ _05414_
+ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__o22ai_4
XANTENNA__12782__B2 _03616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12065__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1235_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08026_ team_01_WB.instance_to_wrap.cpu.K0.code\[2\] _04521_ team_01_WB.instance_to_wrap.cpu.K0.code\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__or3b_4
XFILLER_0_13_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold730 _02078_ vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold741 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout695_A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11337__A2 team_01_WB.instance_to_wrap.cpu.f0.state\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12534__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17956__1456 vssd1 vssd1 vccd1 vccd1 _17956__1456/HI net1456 sky130_fd_sc_hd__conb_1
Xhold752 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[51\] vssd1 vssd1 vccd1 vccd1
+ net2368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold763 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold785 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1402_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold796 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[98\] vssd1 vssd1 vccd1 vccd1
+ net2412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09977_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[2\] net798 net786 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout862_A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08928_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[6\] net911 vssd1
+ vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__and3_1
XANTENNA__13495__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1430 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net3046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[115\] vssd1 vssd1 vccd1 vccd1
+ net3057 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10848__A1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1452 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1463 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08859_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[3\] net911 vssd1
+ vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__and3_1
Xhold1474 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net3090 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16861__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1485 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1496 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3112 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_58_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11870_ net2413 net245 net483 vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13851__C team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08945__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10821_ net529 _07068_ _07159_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11652__B net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11144__S net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13540_ _03926_ _03992_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__xor2_1
X_10752_ _06001_ _06034_ _07091_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ _03930_ _03931_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10683_ net540 _07022_ net549 vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15210_ net1272 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__inv_2
X_12422_ net2239 net293 net420 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__mux2_1
XANTENNA__09769__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16190_ clknet_leaf_115_wb_clk_i _01950_ _00178_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12773__A1 _07251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08680__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12353_ net2115 net305 net430 vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__mux2_1
X_15141_ net1206 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17367__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11304_ _07642_ _07643_ vssd1 vssd1 vccd1 vccd1 _07644_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15072_ net1242 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12284_ net2173 net300 net438 vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14023_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[34\] _04221_ _04233_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[66\]
+ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__a22o_1
X_11235_ net370 _07348_ _07349_ net337 net328 vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12703__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10536__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ net556 _07499_ _07505_ _07071_ vssd1 vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_8_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10117_ _06445_ _06448_ _06453_ _06456_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__or4_1
X_15974_ net1393 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__inv_2
X_11097_ _06901_ _06913_ _07436_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_69_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12828__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10450__C net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17713_ clknet_leaf_82_wb_clk_i _03397_ _01654_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14925_ net1221 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
X_10048_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[0\] net807 net772 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09016__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11500__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold90 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[13\] vssd1 vssd1 vccd1 vccd1
+ net1706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17644_ clknet_leaf_113_wb_clk_i _03329_ _01585_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.bit30
+ sky130_fd_sc_hd__dfrtp_4
X_14856_ net1289 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08855__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13807_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[0\] net833 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[0\] sky130_fd_sc_hd__and2_1
X_17575_ clknet_leaf_77_wb_clk_i _03262_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14787_ net1306 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__inv_2
X_11999_ net2607 net210 net469 vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__mux2_1
XANTENNA__11264__A1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16526_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[24\]
+ _00509_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13738_ net1161 net1162 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.next_lcd_en
+ sky130_fd_sc_hd__and2_1
XFILLER_0_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11989__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16457_ clknet_leaf_133_wb_clk_i _02211_ _00440_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13669_ net1167 _03735_ _04099_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15408_ net1271 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__inv_2
X_16388_ clknet_leaf_77_wb_clk_i net3093 _00371_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12764__A1 _07621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15339_ net1300 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18058_ net1558 vssd1 vssd1 vccd1 vccd1 la_data_out[100] sky130_fd_sc_hd__buf_2
XANTENNA__16734__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _06236_ _06237_ _06238_ _06239_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__or4_1
X_17009_ clknet_leaf_18_wb_clk_i _02696_ _00992_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12613__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10527__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09393__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09831_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[13\] net791 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__a22o_1
Xfanout517 net522 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__clkbuf_4
Xfanout528 net530 vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout539 net540 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_4
X_09762_ _06002_ _06036_ _06068_ _06101_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__or4_1
X_08713_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[5\] net894 vssd1
+ vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09693_ _05657_ _05732_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__xnor2_1
X_08644_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[10\] net892
+ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_29_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08575_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[19\] net934 vssd1
+ vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__and3_1
XANTENNA__10369__A _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout443_A _07959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10058__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09999__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08120__B2 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11899__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16264__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1352_A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout708_A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire918 _04775_ vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire929 _04765_ vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__buf_1
XFILLER_0_17_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13399__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09596__C net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09127_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[14\] net910
+ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__and3_1
XANTENNA_hold1460_A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10766__A0 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_105_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09893__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09058_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[12\] net937
+ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08009_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1 _04506_
+ sky130_fd_sc_hd__inv_2
XANTENNA__12523__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold571 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 net2198
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ _05529_ net372 vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__nor2_1
Xhold593 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08302__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_10__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11366__C net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10270__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__B _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12971_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[115\] net1911 net865 vssd1 vssd1
+ vccd1 vccd1 _02154_ sky130_fd_sc_hd__mux2_1
Xhold1260 _02056_ vssd1 vssd1 vccd1 vccd1 net2876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14710_ net1305 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__inv_2
Xhold1271 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2887 sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ net2864 net321 net482 vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__mux2_1
Xhold1282 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1293 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[78\] vssd1 vssd1 vccd1 vccd1
+ net2909 sky130_fd_sc_hd__dlygate4sd3_1
X_15690_ net1279 vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09133__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08675__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ net1312 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__inv_2
X_11853_ net2549 net296 net490 vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09439__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10279__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10049__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17360_ clknet_leaf_13_wb_clk_i _03047_ _01343_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10804_ _06919_ _07143_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__nor2_1
XANTENNA__11246__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14572_ net1393 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__inv_2
X_11784_ net2259 net298 net497 vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08972__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16311_ clknet_leaf_65_wb_clk_i net2716 _00294_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_13523_ net185 _03977_ _03978_ net725 vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17291_ clknet_leaf_5_wb_clk_i _02978_ _01274_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10735_ _05781_ net332 _07073_ net335 net370 vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__a221o_1
XANTENNA__09787__B net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08662__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16242_ clknet_leaf_80_wb_clk_i net1768 _00230_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
X_10666_ net551 _06313_ _07005_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__o21ba_1
X_13454_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] _05495_ vssd1 vssd1
+ vccd1 vccd1 _03915_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12405_ net2009 net268 net420 vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__mux2_1
X_16173_ clknet_leaf_108_wb_clk_i _01933_ _00161_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13385_ _03845_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__inv_2
X_10597_ net375 _06158_ net544 vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10445__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10221__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15124_ net1264 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__inv_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
X_12336_ net3217 net272 net429 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12941__B net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15055_ net1214 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__inv_2
X_12267_ net2372 net205 net435 vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__mux2_1
XANTENNA__12433__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14214__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14006_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[81\] _04251_ _04260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[57\]
+ _04296_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__a221o_1
XANTENNA__09375__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ _06779_ net335 net332 vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__a21o_1
X_18026__1526 vssd1 vssd1 vccd1 vccd1 _18026__1526/HI net1526 sky130_fd_sc_hd__conb_1
X_12198_ net2577 net274 net445 vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__mux2_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
XANTENNA__11721__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11149_ _07482_ _07486_ _07488_ vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__or3_4
XFILLER_0_78_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14120__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15957_ net1411 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11573__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14908_ net1174 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__inv_2
XANTENNA__10288__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15888_ net1330 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08585__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17627_ clknet_leaf_111_wb_clk_i _03312_ _01568_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_14839_ net1195 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16287__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09978__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17532__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08360_ _04696_ _04697_ _04698_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__or4_1
X_17955__1455 vssd1 vssd1 vccd1 vccd1 _17955__1455/HI net1455 sky130_fd_sc_hd__conb_1
XFILLER_0_54_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17558_ clknet_leaf_139_wb_clk_i _03245_ _01541_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16509_ clknet_leaf_108_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[7\]
+ _00492_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08291_ net1147 net1151 net1153 net1148 vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__nor4b_1
XANTENNA__12608__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17489_ clknet_leaf_17_wb_clk_i _03176_ _01472_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10996__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09850__A1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10917__A _05374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11512__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09189__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10460__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12737__B2 _03585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_6__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10748__B1 _07087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10212__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12343__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13162__B2 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09905__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout303 _07912_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_2
XANTENNA__11467__B net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout314 _07939_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_2
XFILLER_0_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout325 net327 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_2
XANTENNA_fanout393_A _03568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 _06912_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_4
X_09814_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[14\] net808 net793 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__a22o_1
Xfanout347 net348 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_4
Xfanout358 net360 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_2
XANTENNA__09381__A3 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1100_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout369 _06915_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14111__B1 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[20\] net741 _06071_ _06077_
+ _06081_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout560_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08877__C1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[22\] net775 net735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__a22o_1
X_08627_ _04952_ _04963_ _04964_ _04966_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__or4_1
XFILLER_0_51_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09888__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08558_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[19\] net922 vssd1
+ vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10987__A0 _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12518__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08489_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[23\] net691 _04777_ _04792_
+ _04764_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10520_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[31\] net688 net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10451_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[26\] net946
+ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__and3b_1
XFILLER_0_116_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10265__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13170_ net136 net849 net841 net1627 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10382_ net989 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[16\] net941 vssd1
+ vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12121_ net2467 net319 net458 vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12253__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09357__B1 _04806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ net2270 net297 net464 vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__mux2_1
XANTENNA__17405__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold390 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11003_ _05758_ net504 vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__nor2_1
X_16860_ clknet_leaf_37_wb_clk_i _02547_ _00843_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_73_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout870 net871 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_2
XANTENNA__14102__B1 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15811_ net1310 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__inv_2
Xfanout881 net882 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16791_ clknet_leaf_138_wb_clk_i _02478_ _00774_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout892 net893 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15742_ net1274 vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12954_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[5\] _05074_ net1035 vssd1
+ vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__mux2_1
XANTENNA__08178__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2706 sky130_fd_sc_hd__dlygate4sd3_1
X_11905_ net2175 net241 net479 vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__mux2_1
X_15673_ net1259 vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__inv_2
X_12885_ net1859 net870 net357 _03664_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a22o_1
XANTENNA__13208__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08883__A2 _05219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17412_ clknet_leaf_53_wb_clk_i _03099_ _01395_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14624_ net1361 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__inv_2
X_11836_ net2804 net202 net487 vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17343_ clknet_leaf_24_wb_clk_i _03030_ _01326_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14555_ net1408 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__inv_2
XANTENNA__10978__A0 _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ net1991 net206 net495 vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__mux2_1
XANTENNA__12428__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11332__S _07655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14209__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13506_ net198 net194 _07830_ net644 vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__o211a_1
X_17274_ clknet_leaf_60_wb_clk_i _02961_ _01257_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10718_ _06998_ _07002_ net533 vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14486_ net1329 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11698_ net612 _07807_ _07895_ _07894_ vssd1 vssd1 vccd1 vccd1 _07896_ sky130_fd_sc_hd__a31o_2
XFILLER_0_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16225_ clknet_leaf_104_wb_clk_i net1620 _00213_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13437_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\]
+ net597 _03886_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a31oi_1
X_10649_ net511 net510 net543 vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16156_ clknet_leaf_101_wb_clk_i _01919_ _00144_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13368_ net1946 net827 _07650_ _03836_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15107_ net1174 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__inv_2
X_12319_ net2221 net311 net432 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__mux2_1
XANTENNA__12163__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16087_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[9\]
+ _00075_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[9\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10472__A _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13299_ _04516_ _03745_ _03782_ team_01_WB.instance_to_wrap.cpu.f0.next_write_i vssd1
+ vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__o31a_1
XFILLER_0_48_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09348__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17085__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15038_ net1271 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16989_ clknet_leaf_21_wb_clk_i _02676_ _00972_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09530_ net513 _05868_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09461_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[29\] net654 _05795_
+ _05799_ _05800_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09204__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08874__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08412_ _04708_ net729 net720 vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__or3_4
X_09392_ _05570_ _05620_ net559 vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12958__A1 _05219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08343_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[30\] net957 vssd1
+ vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09501__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08626__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12338__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout239_A _07870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08274_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\] net1748 net1047 vssd1 vssd1
+ vccd1 vccd1 _03413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08117__A team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_116_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1050_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_A _03565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16302__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17428__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11394__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_70_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12073__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09339__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout775_A _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1109 net1110 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout188 _07639_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_2
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07989_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1 _04487_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11449__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09728_ net508 _06066_ _06067_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__and3b_1
XFILLER_0_69_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ net510 _05998_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12670_ net2905 net264 net387 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11621_ _07832_ _07834_ net611 vssd1 vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__mux2_4
XANTENNA__12248__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_120_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_18025__1525 vssd1 vssd1 vccd1 vccd1 _18025__1525/HI net1525 sky130_fd_sc_hd__conb_1
XANTENNA__08617__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10557__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10424__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14340_ net1371 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11552_ net1986 net1160 net589 vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10975__A3 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10503_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[31\] net818 net780 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__a22o_1
X_11483_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[21\] net579 vssd1 vssd1 vccd1
+ vccd1 _07769_ sky130_fd_sc_hd__nand2_1
X_14271_ net1376 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16010_ net1396 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__inv_2
X_10434_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\] net777 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__a22o_1
X_13222_ net3134 net353 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1
+ vccd1 vccd1 _01928_ sky130_fd_sc_hd__a22o_1
XANTENNA_input71_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13374__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13079__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13153_ net2029 net844 net839 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[23\] vssd1
+ vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10365_ net768 _06697_ _06701_ _06704_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__nor4_1
XFILLER_0_42_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12104_ net1985 net242 net455 vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__mux2_1
X_17961_ net1461 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
X_13084_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] net2612 net858 vssd1 vssd1
+ vccd1 vccd1 _02041_ sky130_fd_sc_hd__mux2_1
X_10296_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] net626 _06634_ _06635_
+ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__a22o_2
X_17954__1454 vssd1 vssd1 vccd1 vccd1 _17954__1454/HI net1454 sky130_fd_sc_hd__conb_1
XANTENNA__11137__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08538__D1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16912_ clknet_leaf_126_wb_clk_i _02599_ _00895_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12035_ net2955 net204 net464 vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__mux2_1
XANTENNA__11328__A_N team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11688__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17892_ net1595 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XANTENNA__12711__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_69_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09750__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16843_ clknet_leaf_144_wb_clk_i _02530_ _00826_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16945__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11327__S _07655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16774_ clknet_leaf_39_wb_clk_i _02461_ _00757_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13986_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[8\] _04253_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[104\]
+ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__a22o_1
X_15725_ net1221 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12937_ _04968_ _07756_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__nand2_1
XANTENNA__08856__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13849__A_N net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12947__A team_01_WB.instance_to_wrap.cpu.f0.write_data\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15656_ net1289 vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12868_ _04753_ _04944_ _07630_ net578 _03652_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__o311a_1
XFILLER_0_29_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14607_ net1402 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__inv_2
XANTENNA__08863__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11819_ net2907 net310 net493 vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12158__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15587_ net1186 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12799_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] net1056 net365 _03627_
+ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17326_ clknet_leaf_3_wb_clk_i _03013_ _01309_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14538_ net1394 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11997__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17257_ clknet_leaf_23_wb_clk_i _02944_ _01240_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14469_ net1398 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16208_ clknet_leaf_62_wb_clk_i net1812 _00196_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17188_ clknet_leaf_53_wb_clk_i _02875_ _01171_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09033__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11298__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16475__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16139_ clknet_leaf_96_wb_clk_i _01902_ _00127_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17720__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08961_ net603 _05300_ _05266_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13379__A_N team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08892_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[2\] net937 vssd1
+ vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_55_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11745__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08400__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14093__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09513_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[29\] net758 net737 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11300__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout356_A _03741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[29\] net880
+ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09231__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13589__D1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10377__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09375_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[26\] _04778_ net678 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__a22o_1
XANTENNA__12068__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout523_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1265_A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08326_ net1131 net943 vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12800__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17250__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09272__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08257_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[24\] net2007 net1046 vssd1 vssd1
+ vccd1 vccd1 _03430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16818__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08188_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[93\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[85\]
+ net1039 vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09024__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10824__B net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout892_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_103_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09980__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[11\] net795 _06487_ _06488_
+ _06489_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_30_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16968__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13659__A2 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12531__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10081_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[7\] net799 net735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__a22o_1
XANTENNA__08948__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13840_ net1166 net1060 net2066 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[1\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_138_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14084__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13870__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13771_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] _04152_ _04157_ net1170
+ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__o211a_1
X_10983_ _07316_ _07322_ _07310_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__or3b_4
XFILLER_0_74_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15510_ net1247 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12722_ net1156 _04718_ team_01_WB.instance_to_wrap.cpu.DM0.enable team_01_WB.instance_to_wrap.cpu.DM0.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_84_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16490_ clknet_leaf_104_wb_clk_i _02244_ _00473_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16348__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08683__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15441_ net1288 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__inv_2
X_12653_ net2086 net293 net392 vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14982__A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09799__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11604_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\]
+ _07820_ vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__and3_1
XANTENNA__13595__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15372_ net1209 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12584_ net2757 net307 net402 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_142_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09263__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17111_ clknet_leaf_137_wb_clk_i _02798_ _01094_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14323_ net1357 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11070__A2 _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18091_ net636 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_1
XANTENNA__16498__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11535_ net3139 net1157 net587 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] vssd1
+ vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__a22o_1
XANTENNA__12706__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17743__CLK clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17042_ clknet_leaf_134_wb_clk_i _02729_ _01025_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14254_ net1354 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__inv_2
X_11466_ net368 _07760_ net2057 net875 vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_78_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13205_ net3 net837 net630 net2152 vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10417_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[27\] net952
+ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__and3_1
X_14185_ net2904 _04453_ _04455_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11397_ _07668_ _07696_ _07714_ net1062 vssd1 vssd1 vccd1 vccd1 _07722_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10453__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08774__A1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13136_ net104 net847 net633 net1728 vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10348_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[17\] net973
+ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__and3_1
XANTENNA__09019__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12441__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13067_ net2501 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[27\] net864 vssd1 vssd1
+ vccd1 vccd1 _02058_ sky130_fd_sc_hd__mux2_1
X_10279_ net1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[19\] net966
+ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__and3_1
X_17944_ net1444 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
X_12018_ net2974 net300 net470 vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__mux2_1
XANTENNA__08858__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17875_ clknet_leaf_92_wb_clk_i _03550_ _01815_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11530__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16826_ clknet_leaf_45_wb_clk_i _02513_ _00809_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09035__B _05374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11284__C _07621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14075__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16757_ clknet_leaf_126_wb_clk_i _02444_ _00740_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13969_ _04218_ _04224_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__nor2_4
XFILLER_0_92_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11581__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10097__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15708_ net1173 vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11294__C1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16688_ clknet_leaf_127_wb_clk_i _02375_ _00671_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09051__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ net1199 vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_135_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09160_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[16\] net936 vssd1
+ vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_44_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08890__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08057__A3 _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09254__A2 _05591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08111_ net1064 team_01_WB.instance_to_wrap.cpu.f0.num\[8\] vssd1 vssd1 vccd1 vccd1
+ _04581_ sky130_fd_sc_hd__and2_1
X_17309_ clknet_leaf_49_wb_clk_i _02996_ _01292_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09091_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[13\] net938
+ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12616__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10925__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08042_ net1689 net570 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1
+ vccd1 vccd1 _03549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold901 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[94\] vssd1 vssd1 vccd1 vccd1
+ net2517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap620 _04730_ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold923 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold934 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09411__C1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold945 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10021__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold956 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold967 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[35\] vssd1 vssd1 vccd1 vccd1
+ net2583 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09962__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold978 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold989 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _06320_ _06324_ _06329_ _06332_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15228__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08944_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[6\] net927 vssd1
+ vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__and3_1
XANTENNA__12351__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1013_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18024__1524 vssd1 vssd1 vccd1 vccd1 _18024__1524/HI net1524 sky130_fd_sc_hd__conb_1
XFILLER_0_23_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1601 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3217 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09714__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1612 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3228 sky130_fd_sc_hd__dlygate4sd3_1
X_08875_ _05209_ _05210_ _05213_ _05214_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__or4_1
Xhold1623 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3239 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout473_A _07952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1634 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[63\] vssd1 vssd1 vccd1 vccd1
+ net3250 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09190__A1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1645 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net3261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1667 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 net3283
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout640_A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1382_A net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09599__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08150__C1 _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[28\] net695 net678 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[28\]
+ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__a221o_1
X_17953__1453 vssd1 vssd1 vccd1 vccd1 _17953__1453/HI net1453 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_118_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13577__A1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09358_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[25\] net667 net707 vssd1
+ vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08309_ net1131 net962 vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__and2_2
XFILLER_0_62_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12526__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09289_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[22\] net919 vssd1
+ vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11320_ _07656_ net1748 _07655_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11251_ net337 _07351_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10012__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10273__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10202_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[8\] net962 vssd1
+ vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__and3_1
XANTENNA__09953__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11182_ _05006_ _06924_ _07376_ _06919_ _06915_ vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_73_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13865__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10133_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[11\] net951
+ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__and3_1
XANTENNA__12261__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15990_ net1390 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__inv_2
XANTENNA__13501__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08678__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09136__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ _06402_ _06403_ _06343_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__a21o_1
XANTENNA_input34_A gpio_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14941_ net1262 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17660_ clknet_leaf_90_wb_clk_i _03345_ _01601_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14872_ net1176 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17296__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16611_ clknet_leaf_21_wb_clk_i _02298_ _00594_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13823_ net2338 net831 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[16\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_67_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17591_ clknet_leaf_80_wb_clk_i _03278_ _01550_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16542_ clknet_leaf_112_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[8\]
+ _00525_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13754_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__or4b_1
XANTENNA__08186__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10966_ _06314_ _06921_ _07107_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09484__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10729__B _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12705_ net2085 net259 net384 vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16473_ clknet_leaf_81_wb_clk_i _02227_ _00456_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13685_ team_01_WB.instance_to_wrap.cpu.c0.count\[12\] _04107_ vssd1 vssd1 vccd1
+ vccd1 _04108_ sky130_fd_sc_hd__and2_1
XANTENNA__09302__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10897_ net517 _06969_ _06970_ _07236_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15601__A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10448__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15424_ net1242 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13568__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12636_ net2048 net267 net391 vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09236__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12944__B net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15355_ net1181 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__inv_2
X_12567_ net3248 net272 net401 vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__mux2_1
XANTENNA__12436__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14306_ net1353 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__inv_2
X_11518_ net1646 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] team_01_WB.instance_to_wrap.cpu.DM0.next_enable
+ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__mux2_1
X_18074_ net1574 vssd1 vssd1 vccd1 vccd1 la_data_out[116] sky130_fd_sc_hd__buf_2
XANTENNA__12791__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15286_ net1202 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__inv_2
X_12498_ net2544 net206 net407 vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__mux2_1
Xhold208 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[3\] vssd1 vssd1 vccd1 vccd1
+ net1824 sky130_fd_sc_hd__dlygate4sd3_1
X_17025_ clknet_leaf_43_wb_clk_i _02712_ _01008_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold219 net116 vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ net1364 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__inv_2
X_11449_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\] _07672_ net326 vssd1 vssd1 vccd1
+ vccd1 _07749_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14168_ _04189_ _04193_ net1936 vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_128_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ net2017 net844 net631 net1970 vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10480__A _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12171__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[85\] _04245_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[125\]
+ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16513__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ net1615 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
XANTENNA__17639__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18107__1591 vssd1 vssd1 vccd1 vccd1 _18107__1591/HI net1591 sky130_fd_sc_hd__conb_1
XFILLER_0_94_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1270 net1273 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__buf_4
Xfanout1281 net1286 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__buf_2
X_08660_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[10\] net675 _04981_
+ _04983_ _04987_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a2111o_1
Xfanout1292 net1293 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__buf_4
X_17858_ clknet_leaf_83_wb_clk_i team_01_WB.instance_to_wrap.cpu.f0.next_lcd_en _01798_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.enable sky130_fd_sc_hd__dfrtp_1
XANTENNA__14048__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16809_ clknet_leaf_14_wb_clk_i _02496_ _00792_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08591_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[15\] net683 _04928_
+ _04929_ _04930_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_72_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17789_ clknet_leaf_72_wb_clk_i _03465_ _01729_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11515__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10639__B _06928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09212__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08109__B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13559__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09212_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[17\] net886 vssd1
+ vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__and3_1
XANTENNA__17019__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_62_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09143_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[14\] net667 _05457_
+ _05469_ _05477_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_96_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12346__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout221_A _07831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout319_A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09074_ _05405_ _05406_ _05412_ _05413_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_92_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16043__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08025_ team_01_WB.instance_to_wrap.cpu.K0.code\[1\] team_01_WB.instance_to_wrap.cpu.K0.code\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__nand2_1
XANTENNA__17169__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold720 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1130_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[1\] vssd1 vssd1 vccd1 vccd1 net2358
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1228_A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09935__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold753 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold764 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09882__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 net79 vssd1 vssd1 vccd1 vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A _04776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12081__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09976_ _06313_ _06315_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_71_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16193__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08927_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[6\] net883 vssd1
+ vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__and3_1
Xhold1420 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1
+ net3036 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1431 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net3047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1442 _02146_ vssd1 vssd1 vccd1 vccd1 net3058 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08858_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[3\] net927 vssd1
+ vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__and3_1
Xhold1453 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net3069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1464 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1475 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net3091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1486 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[28\] vssd1 vssd1 vccd1 vccd1 net3102
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1497 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[15\] vssd1 vssd1 vccd1 vccd1
+ net3113 sky130_fd_sc_hd__dlygate4sd3_1
X_08789_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[0\] net920 vssd1
+ vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10820_ _06967_ _07159_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_98_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10751_ _06101_ _07089_ _06036_ _06068_ vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__a211oi_2
XANTENNA__09122__C _04799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13470_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _05592_ vssd1 vssd1
+ vccd1 vccd1 _03931_ sky130_fd_sc_hd__or2_1
XANTENNA__09218__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10682_ _04706_ net513 net549 vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12421_ net2397 net315 net421 vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10565__A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12256__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10233__B1 _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15140_ net1237 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12352_ net2140 net309 net428 vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11303_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _05116_ vssd1 vssd1 vccd1
+ vccd1 _07643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15071_ net1254 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12283_ net2381 net279 net436 vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14022_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[90\] _04240_ _04241_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[90\]
+ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11234_ _04738_ _05932_ _06917_ _05707_ _04736_ vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__13087__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11165_ _06905_ _07254_ _07504_ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_8_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[6\] net737 _06454_ _06455_
+ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__a211o_1
X_15973_ net1407 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__inv_2
X_11096_ _07364_ _07379_ _07435_ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_69_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16686__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10047_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[0\] net761 _06380_ _06382_
+ net769 vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__a2111o_1
X_17712_ clknet_leaf_81_wb_clk_i _03396_ _01653_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14924_ net1180 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold80 team_01_WB.instance_to_wrap.cpu.c0.count\[0\] vssd1 vssd1 vccd1 vccd1 net1696
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 net122 vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14855_ net1299 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17643_ clknet_leaf_113_wb_clk_i _03328_ _01584_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_72_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13806_ team_01_WB.EN_VAL_REG net636 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__or2_1
X_17574_ clknet_leaf_60_wb_clk_i _03261_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14786_ net1312 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11998_ net2257 net249 net469 vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__mux2_1
XANTENNA__09457__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16525_ clknet_leaf_116_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[23\]
+ _00508_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13737_ _04511_ _07649_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__or2_1
X_10949_ net330 _07288_ _07287_ _07279_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16456_ clknet_leaf_144_wb_clk_i _02210_ _00439_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13668_ team_01_WB.instance_to_wrap.a1.curr_state\[0\] _03732_ _04098_ vssd1 vssd1
+ vccd1 vccd1 _04099_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_22_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18023__1523 vssd1 vssd1 vccd1 vccd1 _18023__1523/HI net1523 sky130_fd_sc_hd__conb_1
X_15407_ net1218 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12619_ net2325 net315 net398 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__mux2_1
X_16387_ clknet_leaf_85_wb_clk_i net2689 _00370_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12166__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10475__A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13599_ _03907_ _04041_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10224__B1 _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15338_ net1278 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18057_ net1557 vssd1 vssd1 vccd1 vccd1 la_data_out[99] sky130_fd_sc_hd__buf_2
XFILLER_0_124_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15269_ net1207 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17008_ clknet_leaf_127_wb_clk_i _02695_ _00991_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09917__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09393__A1 _05570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09830_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[13\] net790 _06168_
+ _06169_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_6_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout507 _06098_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_4
Xfanout518 net522 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__clkbuf_2
Xfanout529 net530 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17952__1452 vssd1 vssd1 vccd1 vccd1 _17952__1452/HI net1452 sky130_fd_sc_hd__conb_1
XFILLER_0_10_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09761_ _06069_ _06100_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__and2b_1
XANTENNA__09207__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08712_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[5\] net899 vssd1
+ vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__and3_1
XANTENNA__15506__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09692_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] net626 _06030_ _06031_
+ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__a22o_1
XANTENNA__13492__A3 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09504__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[10\] net920 vssd1
+ vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout269_A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08574_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[19\] net907 vssd1
+ vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__and3_1
XANTENNA__09448__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10369__B _05379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16409__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1080_A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout436_A _07963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1178_A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10463__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08781__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12076__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout603_A _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1345_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09126_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[14\] net899
+ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__and3_1
XANTENNA__16559__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09620__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09057_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[12\] net924 vssd1
+ vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08008_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] vssd1 vssd1 vccd1 vccd1 _04505_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_130_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold550 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold583 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09959_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[3\] net789 net776 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__a22o_1
XANTENNA__09117__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12970_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[116\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[124\]
+ net858 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1250 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2866 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09687__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1261 team_01_WB.instance_to_wrap.cpu.f0.num\[21\] vssd1 vssd1 vccd1 vccd1 net2877
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11921_ net1938 net306 net482 vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__mux2_1
Xhold1272 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1283 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1294 _03484_ vssd1 vssd1 vccd1 vccd1 net2910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14640_ net1280 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__inv_2
X_11852_ net3104 net299 net490 vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09439__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _05657_ net509 vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14571_ net1411 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__inv_2
X_11783_ net1863 net281 net496 vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16310_ clknet_leaf_68_wb_clk_i net3173 _00293_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17334__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13522_ net197 net193 _07841_ net643 vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_1195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17290_ clknet_leaf_10_wb_clk_i _02977_ _01273_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10734_ net336 _07073_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__nor2_1
X_16241_ clknet_leaf_81_wb_clk_i net2477 _00229_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13453_ _03900_ _03909_ _03913_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_119_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10665_ net546 _06280_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_58_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12746__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12404_ net2493 net236 net419 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__mux2_1
X_16172_ clknet_leaf_107_wb_clk_i _01932_ _00160_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13384_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _05757_ vssd1 vssd1
+ vccd1 vccd1 _03845_ sky130_fd_sc_hd__or2_1
X_10596_ net374 net342 net546 vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09611__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10757__A1 _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15123_ net1234 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12335_ net2426 net246 net427 vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12714__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15054_ net1295 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__inv_2
X_12266_ net2468 net276 net437 vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__mux2_1
XANTENNA__11706__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14005_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[33\] _04221_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[105\]
+ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__a22o_1
XANTENNA__13171__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11217_ _06814_ _06821_ _07555_ vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12197_ net2695 net209 net445 vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__mux2_1
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
XANTENNA__11182__B2 _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
X_11148_ net330 _07485_ _07487_ _07478_ vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15956_ net1387 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__inv_2
X_11079_ net509 _07095_ _05657_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__and3b_1
XANTENNA__09678__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08866__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11573__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14907_ net1181 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
X_15887_ net1399 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08350__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17626_ clknet_leaf_110_wb_clk_i _03311_ _01567_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14838_ net1201 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14769_ net1324 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__inv_2
X_17557_ clknet_leaf_124_wb_clk_i _03244_ _01540_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16508_ clknet_leaf_108_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[6\]
+ _00491_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08290_ net990 net979 vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17488_ clknet_leaf_15_wb_clk_i _03175_ _01471_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09697__C net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__A1 _06398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16701__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17827__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16439_ clknet_leaf_45_wb_clk_i _02193_ _00422_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12737__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10748__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18109_ net1592 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XANTENNA__12624__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10652__B net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13162__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout304 _07912_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__buf_2
Xfanout315 _07939_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout326 net327 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_2
X_09813_ _06138_ _06150_ _06151_ _06152_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__or4_1
Xfanout337 _06911_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17207__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout348 _04526_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout359 net360 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_4
XANTENNA__10920__A1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10920__B2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[20\] net822 net758 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08877__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09675_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[22\] net953 vssd1
+ vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout553_A _05115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16231__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1295_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17357__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08626_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[11\] net698 net672 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[11\]
+ _04965_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08557_ net1071 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[19\] net886
+ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout720_A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13622__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout818_A _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08488_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[23\] net679 _04818_
+ _04761_ _04786_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09841__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10450_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[26\] net974 vssd1
+ vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__and3b_1
XFILLER_0_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09109_ _05445_ _05446_ _05447_ _05448_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__or4_2
XFILLER_0_116_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10381_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[16\] net785 _06719_
+ _06720_ vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__a211o_1
XANTENNA__12534__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12120_ net2823 net305 net458 vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12051_ net3177 net301 net465 vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__mux2_1
XANTENNA__13153__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold380 _03526_ vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11164__A1 _05262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold391 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[16\] vssd1 vssd1 vccd1 vccd1
+ net2007 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11164__B2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11002_ _05758_ net504 vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18099__1588 vssd1 vssd1 vccd1 vccd1 _18099__1588/HI net1588 sky130_fd_sc_hd__conb_1
Xfanout860 net863 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__clkbuf_4
Xfanout871 net873 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_2
X_15810_ net1310 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__inv_2
XANTENNA__08580__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18022__1522 vssd1 vssd1 vccd1 vccd1 _18022__1522/HI net1522 sky130_fd_sc_hd__conb_1
X_16790_ clknet_leaf_139_wb_clk_i _02477_ _00773_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout882 net883 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__buf_4
XFILLER_0_99_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout893 net894 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__buf_4
XFILLER_0_137_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15741_ net1252 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__inv_2
XANTENNA__08686__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ net1627 net872 net359 _03711_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a22o_1
XANTENNA__08868__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2707 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ net3220 net271 net480 vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_42_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15672_ net1185 vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12884_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[27\] _03663_ net1030 vssd1
+ vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__mux2_1
XANTENNA__08983__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17411_ clknet_leaf_21_wb_clk_i _03098_ _01394_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14623_ net1366 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11835_ net3119 net206 net487 vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__mux2_1
XANTENNA__12709__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output103_A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17342_ clknet_leaf_48_wb_clk_i _03029_ _01325_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10427__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14554_ net1388 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11766_ net3106 net275 net497 vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__mux2_1
XANTENNA__10978__A1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09832__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13505_ _03949_ _03963_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__xnor2_1
X_17273_ clknet_leaf_58_wb_clk_i _02960_ _01256_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17951__1451 vssd1 vssd1 vccd1 vccd1 _17951__1451/HI net1451 sky130_fd_sc_hd__conb_1
X_10717_ _05902_ _06824_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__nand2_1
X_14485_ net1405 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11697_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _07805_ vssd1 vssd1
+ vccd1 vccd1 _07895_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16874__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16224_ clknet_leaf_105_wb_clk_i net1872 _00212_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
X_13436_ _03890_ _03893_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10648_ _06984_ _06987_ net514 vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16155_ clknet_leaf_97_wb_clk_i _01918_ _00143_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12444__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_98_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13367_ net564 team_01_WB.instance_to_wrap.cpu.f0.next_write_i _04486_ vssd1 vssd1
+ vccd1 vccd1 _03836_ sky130_fd_sc_hd__mux2_1
XANTENNA__14225__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10579_ _06910_ _06917_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__or2_4
XFILLER_0_84_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15106_ net1268 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__inv_2
X_12318_ net2552 net294 net431 vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16086_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[8\]
+ _00074_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[8\] sky130_fd_sc_hd__dfrtp_1
X_13298_ net1063 net610 _07710_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15037_ net1263 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__inv_2
X_12249_ net3233 net302 net440 vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09899__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11584__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16988_ clknet_leaf_37_wb_clk_i _02675_ _00971_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09054__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15939_ net1403 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09460_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[29\] _04778_ net669 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[29\]
+ _05783_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08411_ net1156 _04718_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__nor2_2
X_17609_ clknet_leaf_77_wb_clk_i _03296_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12407__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09391_ net559 _05570_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__nor2_1
XANTENNA__12619__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10928__A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08342_ net989 net957 vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__and2_2
XFILLER_0_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1054 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08273_ net2238 net1815 net1046 vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12354__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout301_A _07921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09339__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1210_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11146__A1 _06920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07972__A team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_61_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09890__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout670_A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14096__B1 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout189 net192 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_2
X_07988_ team_01_WB.instance_to_wrap.cpu.f0.i\[7\] vssd1 vssd1 vccd1 vccd1 _04486_
+ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09727_ net378 _05619_ _05731_ _05595_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout935_A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09658_ _04844_ _05733_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_2_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10121__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ _04751_ _04752_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1
+ vccd1 vccd1 _04949_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12529__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ _05918_ _05920_ _05925_ _05928_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__or4_2
XFILLER_0_132_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16897__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11620_ _07820_ _07833_ vssd1 vssd1 vccd1 vccd1 _07834_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08078__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09814__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10557__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_132_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11551_ net1829 net1160 vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__and2_1
XANTENNA__09130__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10502_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[31\] net746 _06834_ _06838_
+ _06840_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__a2111o_1
X_14270_ net1321 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__inv_2
XANTENNA__14020__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13868__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11482_ net367 _07768_ net2260 net874 vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13221_ net2386 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1
+ vccd1 vccd1 _01929_ sky130_fd_sc_hd__a22o_1
X_10433_ _06769_ _06770_ _06771_ _06772_ vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__or4_1
XANTENNA__13374__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12264__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13152_ net1957 net844 net839 net1886 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__a22o_1
XANTENNA_input64_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10364_ _06691_ _06692_ _06702_ _06703_ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ net3101 net271 net457 vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17960_ net1460 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
X_13083_ net2721 net2681 net864 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10295_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] net764 net622 vssd1
+ vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__o21a_1
XANTENNA__08978__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12034_ net2077 net207 net464 vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__mux2_1
X_16911_ clknet_leaf_141_wb_clk_i _02598_ _00894_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_17891_ net1594 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_109_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11608__S _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08553__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16842_ clknet_leaf_11_wb_clk_i _02529_ _00825_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10360__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout690 _04773_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_8
X_16773_ clknet_leaf_31_wb_clk_i _02460_ _00756_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13985_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[8\] _04226_ _04256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[40\]
+ _04276_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12936_ net359 _03699_ _03700_ net872 net2038 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a32o_1
X_15724_ net1210 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__inv_2
XANTENNA__15604__A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10112__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12947__B net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09602__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15655_ net1327 vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__inv_2
XANTENNA__12439__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12867_ net583 _07756_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11818_ net2523 net297 net494 vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14606_ net1401 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__inv_2
XANTENNA__09266__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15586_ net1267 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12798_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[10\] _07531_ net1033 vssd1 vssd1
+ vccd1 vccd1 _03627_ sky130_fd_sc_hd__mux2_1
XANTENNA__09805__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14537_ net1399 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__inv_2
X_17325_ clknet_leaf_138_wb_clk_i _03012_ _01308_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11749_ _04501_ _07936_ net616 vssd1 vssd1 vccd1 vccd1 _07937_ sky130_fd_sc_hd__mux2_2
XFILLER_0_56_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14468_ net1335 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__inv_2
XANTENNA__17052__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17256_ clknet_leaf_22_wb_clk_i _02943_ _01239_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14011__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16207_ clknet_leaf_62_wb_clk_i net1776 _00195_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
X_13419_ _03877_ _03878_ _03869_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_12_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17187_ clknet_leaf_19_wb_clk_i _02874_ _01170_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12174__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14399_ net1365 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10179__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09049__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16138_ clknet_leaf_94_wb_clk_i _01901_ _00126_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08792__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13117__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08960_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] net705 _05296_ _05299_
+ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__o22a_2
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16069_ clknet_leaf_121_wb_clk_i _01862_ _00057_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_0_110_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13522__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08891_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[2\] net916 vssd1
+ vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11518__S team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14078__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10351__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09512_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[29\] net762 net752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[29\]
+ _05850_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11300__A1 _05153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09443_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[29\] net898
+ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout251_A _07904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12349__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09257__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09374_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[26\] net693 net659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08325_ net1151 net1153 net1146 net1148 vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__and4b_4
XFILLER_0_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout516_A _05261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1160_A team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1258_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08256_ net2353 net2244 net1050 vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14002__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18021__1521 vssd1 vssd1 vccd1 vccd1 _18021__1521/HI net1521 sky130_fd_sc_hd__conb_1
XFILLER_0_132_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09885__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12084__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08187_ net2517 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[86\] net1042 vssd1 vssd1
+ vccd1 vccd1 _03500_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout885_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08798__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10080_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[7\] net969 vssd1
+ vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08535__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17950__1450 vssd1 vssd1 vccd1 vccd1 _17950__1450/HI net1450 sky130_fd_sc_hd__conb_1
XANTENNA__14069__B1 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09125__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13770_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[3\] _04146_ vssd1 vssd1
+ vccd1 vccd1 _04157_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_1228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10982_ net556 _07311_ _07321_ net330 vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08964__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12721_ team_01_WB.instance_to_wrap.a1.WRITE_I team_01_WB.instance_to_wrap.cpu.RU0.state\[1\]
+ _03571_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__or3_1
XFILLER_0_116_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12259__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15440_ net1226 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ net1992 net315 net394 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09248__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11603_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\]
+ _07819_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__and3_1
X_15371_ net1295 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ net2155 net313 net400 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17110_ clknet_leaf_1_wb_clk_i _02797_ _01093_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14322_ net1356 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__inv_2
X_11534_ net1759 net1157 net587 net1141 vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18090_ net637 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17041_ clknet_leaf_13_wb_clk_i _02728_ _01024_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11399__A team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14253_ net1354 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__inv_2
X_11465_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[30\] net580 vssd1 vssd1 vccd1
+ vccd1 _07760_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_78_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13204_ net4 net836 net629 net1798 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__o22a_1
X_10416_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[27\] net963
+ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14184_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\] _04453_ net1410 vssd1
+ vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11396_ _07668_ _07697_ _07699_ _07714_ vssd1 vssd1 vccd1 vccd1 _07721_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_81_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08774__A2 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13135_ net1769 net847 net632 team_01_WB.instance_to_wrap.a1.ADR_I\[8\] vssd1 vssd1
+ vccd1 vccd1 _02006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10347_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[17\] net959
+ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__and3_1
XANTENNA__14503__A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13066_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[20\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[28\]
+ net854 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__mux2_1
X_17943_ net1443 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
X_10278_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[19\] net964
+ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11338__S _07655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12017_ net2205 net280 net467 vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__mux2_1
X_17874_ clknet_leaf_94_wb_clk_i _03549_ _01814_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11530__B2 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16825_ clknet_leaf_47_wb_clk_i _02512_ _00808_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15334__A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16756_ clknet_leaf_128_wb_clk_i _02443_ _00739_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13968_ _04225_ _04232_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__nor2_4
XFILLER_0_57_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17418__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10097__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15707_ net1178 vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12919_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[17\] net1031 vssd1 vssd1 vccd1
+ vccd1 _03689_ sky130_fd_sc_hd__or2_1
XANTENNA__12169__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13899_ net571 _04200_ _04201_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__and3_1
X_16687_ clknet_leaf_142_wb_clk_i _02374_ _00670_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09239__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15638_ net1201 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_135_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15569_ net1292 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16442__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17568__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11801__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08110_ net1064 team_01_WB.instance_to_wrap.cpu.f0.num\[8\] vssd1 vssd1 vccd1 vccd1
+ _04580_ sky130_fd_sc_hd__nor2_1
X_17308_ clknet_leaf_36_wb_clk_i _02995_ _01291_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09090_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[13\] net885 vssd1
+ vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08041_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[14\] net569 net347 net3289
+ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__a22o_1
X_17239_ clknet_leaf_136_wb_clk_i _02926_ _01222_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold902 _03500_ vssd1 vssd1 vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold913 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold924 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold935 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 net2551
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[14\] vssd1 vssd1 vccd1 vccd1
+ net2562 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08765__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold957 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold968 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[2\] net737 _06330_ _06331_
+ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__a211o_1
XANTENNA__12632__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold979 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08943_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[6\] net905 vssd1
+ vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__and3_1
XANTENNA__09507__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout299_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08874_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[3\] net695 net684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[3\]
+ _05204_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__a221o_1
Xhold1602 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1613 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3229 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1006_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1624 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1635 _03477_ vssd1 vssd1 vccd1 vccd1 net3251 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1646 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3262 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09190__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1657 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3273 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1668 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 net3284
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09478__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17098__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12079__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout633_A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1375_A net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09426_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[28\] net900
+ net651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[28\] vssd1 vssd1 vccd1
+ vccd1 _05766_ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13577__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09357_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[25\] net692 _04806_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout800_A _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12785__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ net1148 net1154 net1151 net1146 vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_35_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09288_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[22\] net878 vssd1
+ vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16935__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08239_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[42\] net1667 net1043 vssd1 vssd1
+ vccd1 vccd1 _03448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11250_ _05967_ _06748_ _06749_ vssd1 vssd1 vccd1 vccd1 _07590_ sky130_fd_sc_hd__and3_1
XANTENNA__09402__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10201_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[8\] net969 vssd1
+ vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_73_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11181_ _06532_ _07190_ net345 vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__a21o_1
XANTENNA__12542__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10132_ _06442_ _06471_ _06470_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08321__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10570__B _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10063_ _06339_ _06342_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__xnor2_1
X_14940_ net1173 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__inv_2
XANTENNA__11512__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14871_ net1195 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16610_ clknet_leaf_34_wb_clk_i _02297_ _00593_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15154__A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11682__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13822_ net2326 net834 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[15\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_82_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17590_ clknet_leaf_80_wb_clk_i _03277_ _01549_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13265__A1 _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13265__B2 _04621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13753_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1 _04142_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16541_ clknet_leaf_109_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[7\]
+ _00524_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_10965_ _05263_ _07303_ _07304_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_97_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12704_ net2526 net232 net385 vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__mux2_1
X_16472_ clknet_leaf_83_wb_clk_i _02226_ _00455_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13684_ team_01_WB.instance_to_wrap.cpu.c0.count\[10\] team_01_WB.instance_to_wrap.cpu.c0.count\[11\]
+ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10896_ net517 _07138_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15423_ net1254 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__inv_2
X_12635_ net2714 net235 net391 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__mux2_1
XANTENNA__13568__A2 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12717__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11579__A1 _06961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11621__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13402__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15354_ net1193 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12566_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[21\] net243 net399 vssd1
+ vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09641__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08995__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11517_ net1682 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\] team_01_WB.instance_to_wrap.cpu.DM0.next_enable
+ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__mux2_1
X_14305_ net1357 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__inv_2
X_15285_ net1219 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__inv_2
X_18073_ net1573 vssd1 vssd1 vccd1 vccd1 la_data_out[115] sky130_fd_sc_hd__buf_2
XFILLER_0_13_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12497_ net2951 net274 net409 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17024_ clknet_leaf_33_wb_clk_i _02711_ _01007_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold209 team_01_WB.instance_to_wrap.a1.ADR_I\[23\] vssd1 vssd1 vccd1 vccd1 net1825
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14236_ net1367 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__inv_2
X_11448_ _07674_ _07748_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14167_ _04189_ _04193_ _04444_ net1412 vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12452__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15329__A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10761__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11379_ _07707_ vssd1 vssd1 vccd1 vccd1 _07708_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11751__A1 _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13118_ net1799 net843 net631 team_01_WB.instance_to_wrap.a1.ADR_I\[25\] vssd1 vssd1
+ vccd1 vccd1 _02023_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11576__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14098_ _04378_ _04380_ _04382_ _04384_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_52_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[37\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[45\]
+ net854 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__mux2_1
X_17926_ net1614 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_33_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1260 net1261 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__buf_4
Xfanout1271 net1273 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__buf_2
Xfanout1282 net1286 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__buf_4
X_17857_ clknet_leaf_76_wb_clk_i net1710 _01797_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[127\]
+ sky130_fd_sc_hd__dfrtp_1
X_18020__1520 vssd1 vssd1 vccd1 vccd1 _18020__1520/HI net1520 sky130_fd_sc_hd__conb_1
Xfanout1293 net1294 vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_117_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11592__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16808_ clknet_leaf_31_wb_clk_i _02495_ _00791_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16808__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08590_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[15\] net674 net658 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__a22o_1
X_17788_ clknet_leaf_66_wb_clk_i _03464_ _01728_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09062__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16739_ clknet_leaf_21_wb_clk_i _02426_ _00722_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16958__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09211_ net1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[17\] net894
+ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_27_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12627__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09142_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[14\] net680 _05463_
+ _05465_ _05476_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_96_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09073_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[12\] net676 _05383_
+ _05386_ _05394_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__a2111o_1
XANTENNA__16045__D net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout214_A _07838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08024_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] _04506_ _04511_ _04517_ _04519_
+ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold710 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 net2326
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13192__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold743 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[62\] vssd1 vssd1 vccd1 vccd1
+ net2359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold754 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12362__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1123_A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold765 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold776 _02011_ vssd1 vssd1 vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16338__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold787 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08779__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09975_ net526 _06282_ _06314_ net378 vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold798 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
X_08926_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] net599 net596 vssd1 vssd1
+ vccd1 vccd1 _05266_ sky130_fd_sc_hd__and3_1
XANTENNA__13495__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1410 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1421 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09163__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08857_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[3\] net911 vssd1
+ vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__and3_1
Xhold1432 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3048 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout750_A _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1443 team_01_WB.instance_to_wrap.cpu.f0.num\[25\] vssd1 vssd1 vccd1 vccd1 net3059
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1454 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1465 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[73\] vssd1 vssd1 vccd1 vccd1
+ net3081 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout848_A _03731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08910__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1476 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[103\] vssd1 vssd1 vccd1 vccd1
+ net3092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1487 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3103 sky130_fd_sc_hd__dlygate4sd3_1
X_08788_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[0\] net696 _05125_ _05126_
+ _05127_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_54_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1498 _02054_ vssd1 vssd1 vccd1 vccd1 net3114 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13247__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_79_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10750_ _06101_ _07089_ _06068_ vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09871__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09409_ _05742_ _05744_ _05746_ _05748_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__or4_1
XFILLER_0_133_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17883__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10681_ _05901_ _06825_ _06827_ net344 vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__a31o_1
XANTENNA__12537__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17899__1419 vssd1 vssd1 vccd1 vccd1 _17899__1419/HI net1419 sky130_fd_sc_hd__conb_1
XFILLER_0_30_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12420_ net2288 net318 net421 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09623__B1 _05961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10565__B net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12351_ net2899 net297 net430 vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11430__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_67_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_75_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ _07640_ _07641_ vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__and2b_1
X_15070_ net1251 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__inv_2
X_12282_ net3109 net302 net436 vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14021_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[42\] _04256_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[106\]
+ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__a22o_1
X_11233_ _06966_ _07265_ vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__nand2_1
XANTENNA__11677__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10581__A _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12272__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10536__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12930__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08689__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11164_ _05262_ _07467_ _07503_ net531 vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__a22o_1
XANTENNA__17263__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[6\] net816 net784 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__a22o_1
X_11095_ _07334_ _07391_ _07398_ _07434_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__and4b_1
X_15972_ net1387 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17711_ clknet_leaf_82_wb_clk_i _03395_ _01652_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14923_ net1295 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
X_10046_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[0\] net757 _06370_ _06377_
+ _06381_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_69_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold70 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[88\] vssd1 vssd1 vccd1 vccd1 net1686
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 net1697
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 _01988_ vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ clknet_leaf_111_wb_clk_i _03327_ _01583_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\]
+ sky130_fd_sc_hd__dfrtp_4
X_14854_ net1299 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13238__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_1616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13805_ _04159_ _04181_ _04183_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a21bo_1
X_17573_ clknet_leaf_60_wb_clk_i _03260_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11997_ net2539 net215 net469 vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__mux2_1
X_14785_ net1250 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16524_ clknet_leaf_116_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[22\]
+ _00507_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10948_ _07283_ _07286_ net526 vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__mux2_1
X_13736_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid net3290 _04523_ _04135_ vssd1
+ vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__a31o_1
XANTENNA__09862__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16455_ clknet_leaf_11_wb_clk_i _02209_ _00438_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12447__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10879_ _07028_ _07036_ net517 vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__mux2_1
X_13667_ net3208 _04097_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10756__A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14228__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12749__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15406_ net1285 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12618_ net3122 net320 net398 vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16386_ clknet_leaf_62_wb_clk_i _02140_ _00369_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[109\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_5_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09614__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13598_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _05381_ _04029_ vssd1
+ vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15337_ net1229 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__inv_2
X_12549_ net2336 net294 net406 vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18056_ net1556 vssd1 vssd1 vccd1 vccd1 la_data_out[98] sky130_fd_sc_hd__buf_2
XANTENNA_1 _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15268_ net1239 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__inv_2
XANTENNA__13174__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17007_ clknet_leaf_142_wb_clk_i _02694_ _00990_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15059__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14219_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] vssd1 vssd1 vccd1
+ vccd1 _02268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12182__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10491__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15199_ net1257 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10527__A2 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09057__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout508 _06065_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__buf_2
Xfanout519 net520 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09760_ _06099_ net507 vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_24_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08711_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[5\] net883 vssd1
+ vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__and3_1
XANTENNA__09145__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17909_ net1601 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
X_09691_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] net765 net622 vssd1
+ vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__o21a_1
Xfanout1090 net1092 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08642_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[10\] net935
+ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08573_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[19\] net915 vssd1
+ vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15522__A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout331_A _06924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout429_A _07965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09125_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[14\] net924
+ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1240_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09056_ net1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[12\] net891
+ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__and3_1
XANTENNA__17286__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09893__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout798_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13165__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ net1161 vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12092__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold540 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold551 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11715__A1 _07290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09384__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold573 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold584 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold595 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout965_A _04645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08302__C net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08592__B1 _04808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[3\] net738 _06291_ _06295_
+ _06297_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_99_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08909_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[2\] net669 _05231_ _05235_
+ _05237_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_99_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09889_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[5\] net942 vssd1
+ vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_114_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1240 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[89\] vssd1 vssd1 vccd1 vccd1
+ net2856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[75\] vssd1 vssd1 vccd1 vccd1
+ net2867 sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ net2993 net310 net481 vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__mux2_1
Xhold1262 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2878 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10151__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1273 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1284 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1295 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2911 sky130_fd_sc_hd__dlygate4sd3_1
X_11851_ net2682 net282 net487 vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__mux2_1
XANTENNA__09133__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10279__C net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10802_ _05657_ net509 vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__or2_1
X_14570_ net1388 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11782_ net2109 net303 net496 vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09844__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08972__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13521_ _03944_ _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10733_ _05781_ _05898_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12267__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16240_ clknet_leaf_81_wb_clk_i _02000_ _00228_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
X_13452_ _03904_ _03906_ _03912_ _03911_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__a31oi_1
X_10664_ _07000_ _07003_ net517 vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__mux2_1
XANTENNA__17629__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12403_ net2051 net241 net419 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13383_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] _05780_ vssd1 vssd1
+ vccd1 vccd1 _03844_ sky130_fd_sc_hd__xor2_1
X_16171_ clknet_leaf_90_wb_clk_i net3062 _00159_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10595_ net553 _06902_ vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_88_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10757__A2 _05996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15122_ net1232 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__inv_2
X_12334_ net2292 net202 net427 vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13156__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15053_ net1212 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12265_ net3135 net209 net437 vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__mux2_1
XANTENNA__16653__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10509__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11706__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14004_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[9\] _04253_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12903__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11216_ _06814_ _07555_ _06821_ vssd1 vssd1 vccd1 vccd1 _07556_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09375__A2 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12196_ net1953 net249 net445 vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__mux2_1
XANTENNA__11182__A2 _06924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
X_11147_ _06906_ _07319_ _07483_ net525 vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__o22a_1
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__15607__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14511__A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14120__A2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09605__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15955_ net1403 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__inv_2
X_11078_ _07415_ _07416_ _07417_ _07357_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__o31a_1
X_10029_ _06366_ _06367_ _06368_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__and3_1
XANTENNA__10250__S net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14906_ net1192 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
X_15886_ net1394 vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__inv_2
XANTENNA__10142__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17625_ clknet_leaf_111_wb_clk_i _03310_ _01566_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14837_ net1221 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__inv_2
XANTENNA__09043__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16033__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17159__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12966__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17556_ clknet_leaf_128_wb_clk_i _03243_ _01539_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09835__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14768_ net1274 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__inv_2
XANTENNA__09978__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16507_ clknet_leaf_109_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[5\]
+ _00490_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09340__A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13719_ team_01_WB.instance_to_wrap.cpu.c0.count\[10\] _04106_ net3098 vssd1 vssd1
+ vccd1 vccd1 _04129_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12177__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17487_ clknet_leaf_141_wb_clk_i _03174_ _01470_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14699_ net1318 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10996__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16438_ clknet_leaf_47_wb_clk_i _02192_ _00421_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16183__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16369_ clknet_leaf_56_wb_clk_i _02123_ _00352_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[92\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__12905__S net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18108_ net638 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08810__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13147__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18039_ net1539 vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__buf_2
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout305 _07935_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout316 _07939_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_2
XANTENNA__11173__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10905__C1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09812_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[14\] net823 net798 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__a22o_1
Xfanout327 _07698_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_2
XANTENNA__12640__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout338 _06911_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__buf_2
Xfanout349 _03742_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_2
XFILLER_0_94_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17898__1418 vssd1 vssd1 vccd1 vccd1 _17898__1418/HI net1418 sky130_fd_sc_hd__conb_1
XANTENNA__14111__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[20\] net777 net748 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_129_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12122__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout281_A _07917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[22\] net967 vssd1
+ vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08625_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[11\] net694 net675 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__a22o_1
XANTENNA__10684__A1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1190_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout546_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1288_A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15252__A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08556_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[19\] net915
+ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__and3_1
XANTENNA__08629__A1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13622__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__C net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16526__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11633__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_122_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12087__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08487_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[23\] net694 _04774_ _04781_
+ _04826_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_135_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_138_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12189__A1 _07941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16676__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[13\] net658 _05420_
+ _05426_ _05439_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_33_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10380_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[16\] net784 net747 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13138__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09039_ _05264_ _05265_ _05302_ _05377_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__or4b_4
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12050_ net2006 net281 net463 vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__mux2_1
XANTENNA__09357__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold370 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[1\] vssd1 vssd1 vccd1 vccd1
+ net1986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09128__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold392 _03430_ vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08565__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ _07072_ _07073_ _07340_ _07045_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__o211ai_1
XANTENNA__12550__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout850 net851 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
Xfanout861 net863 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14102__A2 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout872 net873 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__buf_4
Xfanout883 _04803_ vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__buf_4
Xfanout894 _04793_ vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__buf_4
X_15740_ net1175 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__inv_2
XANTENNA__10124__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12952_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[6\] _05300_ net1035 vssd1
+ vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10675__A1 _07014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11903_ net3145 net245 net479 vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__mux2_1
Xhold1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15671_ net1196 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12883_ _05756_ net577 net361 vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_119_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17410_ clknet_leaf_36_wb_clk_i _03097_ _01393_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14622_ net1366 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11834_ net2330 net275 net488 vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13613__A1 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09160__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17341_ clknet_leaf_21_wb_clk_i _03028_ _01324_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14553_ net1399 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__inv_2
X_11765_ net2625 net209 net498 vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_82_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13504_ _03842_ _03843_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__and2_1
X_10716_ _07020_ _07021_ _07053_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__o21ai_4
X_17272_ clknet_leaf_28_wb_clk_i _02959_ _01255_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14484_ net1390 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_11_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11696_ net720 _07520_ net615 _07893_ vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16223_ clknet_leaf_106_wb_clk_i net1836 _00211_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ _06985_ _06986_ net538 vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13435_ _03889_ _03892_ _03895_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__or3_1
XFILLER_0_64_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13410__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16154_ clknet_leaf_99_wb_clk_i _01917_ _00142_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13366_ net1722 _03835_ net826 vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10578_ _06910_ _06917_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__nor2_1
XANTENNA__13129__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15105_ net1250 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__inv_2
X_12317_ net2923 net299 net433 vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16085_ clknet_leaf_102_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[7\]
+ _00073_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[7\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09319__B _05570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13297_ net585 _07649_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.next_write_i
+ sky130_fd_sc_hd__or2_1
XFILLER_0_122_1517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09348__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12248_ net2793 net284 net442 vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__mux2_1
X_15036_ net1173 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12179_ net2504 net253 net449 vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__mux2_1
XANTENNA__12460__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14241__A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10363__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16987_ clknet_leaf_17_wb_clk_i _02674_ _00970_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13301__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15938_ net1390 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10115__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16549__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15869_ net1345 vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11804__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ _04736_ net562 vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__nand2_2
X_17608_ clknet_leaf_72_wb_clk_i _03295_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09390_ net377 net343 _05493_ net559 vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08341_ net1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[30\] net945
+ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__and3_1
X_17539_ clknet_leaf_23_wb_clk_i _03226_ _01522_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09501__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16699__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08272_ net2164 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] net1052 vssd1 vssd1
+ vccd1 vccd1 _03415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13368__B1 _07650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12635__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09587__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10155__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09339__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout496_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13872__A_N net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12370__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1203_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07987_ net1064 vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout663_A _04808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18105__1590 vssd1 vssd1 vccd1 vccd1 _18105__1590/HI net1590 sky130_fd_sc_hd__conb_1
X_09726_ _05570_ _05618_ _05594_ net559 vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__a211o_1
XANTENNA__10106__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09511__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09657_ net510 vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout928_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11714__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__inv_2
X_09588_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[25\] net789 net770 _05926_
+ _05927_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__a2111o_1
X_08539_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[18\] net677 _04856_
+ _04865_ _04870_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08078__A2 team_01_WB.instance_to_wrap.cpu.K0.keyvalid vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11550_ net1824 net1160 vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__and2_1
XANTENNA__11082__A1 _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10501_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[31\] net964
+ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__and3_1
XANTENNA__12545__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11481_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[22\] net579 vssd1 vssd1 vccd1
+ vccd1 _07768_ sky130_fd_sc_hd__nand2_1
XANTENNA__10854__A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14326__A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ net2360 net354 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[30\] vssd1 vssd1
+ vccd1 vccd1 _01930_ sky130_fd_sc_hd__a22o_1
X_10432_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[27\] net792 net780 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08324__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12582__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13151_ net125 net847 net842 net1801 vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__a22o_1
X_10363_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[17\] net785 net746 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12102_ net3198 net243 net455 vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13082_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[12\]
+ net854 vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__mux2_1
X_10294_ _06621_ _06626_ _06633_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__or3_4
XANTENNA_input57_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12033_ net2650 net274 net465 vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__mux2_1
X_16910_ clknet_leaf_3_wb_clk_i _02597_ _00893_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12280__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17890_ net107 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09750__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16841_ clknet_leaf_14_wb_clk_i _02528_ _00824_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout680 _04789_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__buf_8
Xfanout691 _04772_ vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_8
X_16772_ clknet_leaf_52_wb_clk_i _02459_ _00755_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08994__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13984_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[32\] _04230_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[56\]
+ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15723_ net1300 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12935_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[12\] net1036 vssd1 vssd1 vccd1
+ vccd1 _03700_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13405__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15654_ net1325 vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12866_ net1166 team_01_WB.instance_to_wrap.cpu.RU0.state\[6\] team_01_WB.instance_to_wrap.a1.WRITE_I
+ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14605_ net1348 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__inv_2
X_11817_ net2779 net299 net494 vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15585_ net1251 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__inv_2
X_12797_ net1792 net639 net606 _03626_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17324_ clknet_leaf_130_wb_clk_i _03011_ _01307_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14536_ net1384 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[2\] _07489_ net718 vssd1 vssd1
+ vccd1 vccd1 _07936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17897__1417 vssd1 vssd1 vccd1 vccd1 _17897__1417/HI net1417 sky130_fd_sc_hd__conb_1
X_17255_ clknet_leaf_16_wb_clk_i _02942_ _01238_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14467_ net1392 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__inv_2
XANTENNA__12455__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11679_ net2829 net263 net501 vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16206_ clknet_leaf_79_wb_clk_i net2016 _00194_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13418_ _03869_ _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_12_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17186_ clknet_leaf_34_wb_clk_i _02873_ _01169_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14398_ net1338 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16221__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16137_ clknet_leaf_98_wb_clk_i _01900_ _00125_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13349_ net1684 net826 _03822_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16068_ clknet_leaf_118_wb_clk_i _01861_ _00056_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11595__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09726__C1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15019_ net1300 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__inv_2
X_08890_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[2\] net903 vssd1
+ vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16371__CLK clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10887__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08369__A_N team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10004__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09511_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[29\] net738 _05841_
+ _05842_ _05845_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_91_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11300__A2 _05154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[29\] net904
+ net664 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[29\] vssd1 vssd1 vccd1
+ vccd1 _05782_ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09373_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[26\] net668 _05709_ _05710_
+ _05712_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09231__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout244_A _07862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10377__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08324_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[30\] net945 vssd1
+ vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12800__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[26\] net2229 net1043 vssd1 vssd1
+ vccd1 vccd1 _03432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12365__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08186_ net3186 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[87\] net1047 vssd1 vssd1
+ vccd1 vccd1 _03501_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07983__A team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09980__A2 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout780_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16714__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout878_A _04810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11709__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13513__B1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14069__B2 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09709_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[21\] net799 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__a22o_1
X_10981_ _06905_ _07317_ _07320_ vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__a21o_1
XANTENNA__10849__A _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ team_01_WB.instance_to_wrap.cpu.RU0.state\[6\] team_01_WB.instance_to_wrap.cpu.RU0.state\[2\]
+ net1061 net1165 vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_84_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ net2240 net318 net394 vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _07818_ vssd1 vssd1
+ vccd1 vccd1 _07819_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09799__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15370_ net1226 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__inv_2
X_12582_ net2378 net296 net402 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__mux2_1
XANTENNA__09653__D1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14321_ net1356 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11533_ net2018 net1157 net587 net1116 vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__a22o_1
XANTENNA__12275__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire322 _07464_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_48_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14056__A _04226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17040_ clknet_leaf_127_wb_clk_i _02727_ _01023_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11464_ _07754_ net368 net2105 net875 vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__o2bb2a_1
X_14252_ net1352 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_78_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10415_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[27\] net976
+ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__and3_1
X_13203_ net5 net836 net629 net3270 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14183_ _04453_ _04454_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__nor2_1
X_11395_ net325 _07715_ _07720_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__and3_1
XANTENNA__08989__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16394__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13134_ net106 net847 net632 net1795 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a22o_1
X_10346_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[17\] net943
+ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13065_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[21\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[29\]
+ net854 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__mux2_1
X_17942_ net1442 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__10318__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10277_ net1120 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[19\] net971
+ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__and3_1
X_12016_ net2083 net303 net468 vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__mux2_1
X_17873_ clknet_leaf_95_wb_clk_i _03548_ _01813_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11530__A2 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16824_ clknet_leaf_27_wb_clk_i _02511_ _00807_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16755_ clknet_leaf_135_wb_clk_i _02442_ _00738_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13967_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ _04220_ _04223_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__and4_4
XFILLER_0_18_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15706_ net1190 vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__inv_2
XANTENNA__10097__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12918_ net361 _03687_ net1029 vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16686_ clknet_leaf_8_wb_clk_i _02373_ _00669_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13898_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\] _04141_ vssd1 vssd1 vccd1
+ vccd1 _04201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15637_ net1223 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__inv_2
XANTENNA__09051__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12849_ net3243 net266 net379 vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10197__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ net1224 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08890__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17307_ clknet_leaf_50_wb_clk_i _02994_ _01290_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14519_ net1332 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12794__B2 _03624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12185__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10494__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15499_ net1299 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08040_ net1692 net568 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1
+ vccd1 vccd1 _03551_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17238_ clknet_leaf_1_wb_clk_i _02925_ _01221_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16737__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold903 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
X_17169_ clknet_leaf_19_wb_clk_i _02856_ _01152_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold914 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10021__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold947 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold958 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[43\] vssd1 vssd1 vccd1 vccd1
+ net2574 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09962__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09991_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[2\] net754 net748 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold969 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 net2585
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08942_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[6\] net927 vssd1
+ vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_1290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09175__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[3\] net681 _05194_ _05195_
+ _05206_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__a2111o_1
Xhold1603 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1614 team_01_WB.instance_to_wrap.cpu.f0.num\[15\] vssd1 vssd1 vccd1 vccd1 net3230
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1625 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[43\] vssd1 vssd1 vccd1 vccd1
+ net3241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1636 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3252 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15525__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1647 team_01_WB.instance_to_wrap.cpu.f0.write_data\[8\] vssd1 vssd1 vccd1 vccd1
+ net3263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1658 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3274 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1669 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 net3285
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout459_A _07955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09425_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[28\] net672 net662 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[28\]
+ _05762_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__a221o_1
XANTENNA__16267__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout626_A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1368_A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07978__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09356_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[25\] net683 _05694_
+ _05695_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_118_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_139_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_139_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13982__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08307_ net1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[30\] net964
+ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__and3_1
XANTENNA__12095__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09287_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[22\] net897 vssd1
+ vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08238_ net3241 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[35\] net1051 vssd1 vssd1
+ vccd1 vccd1 _03449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17662__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout995_A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08169_ net2531 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[104\] net1052 vssd1 vssd1
+ vccd1 vccd1 _03518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10548__A0 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10200_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[8\] net957 vssd1
+ vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__and3_1
XANTENNA__10012__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11180_ net563 _07173_ _07510_ _07519_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__a31o_2
XFILLER_0_82_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09953__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10131_ net373 _06467_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__nor2_1
XANTENNA__08321__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10062_ _06399_ _06400_ _06369_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__a21o_1
XANTENNA__09136__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14870_ net1197 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
X_17896__1416 vssd1 vssd1 vccd1 vccd1 _17896__1416/HI net1416 sky130_fd_sc_hd__conb_1
XFILLER_0_118_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17042__CLK clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13821_ net2343 net833 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[14\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__11682__B _07809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16540_ clknet_leaf_108_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[6\]
+ _00523_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_67_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13752_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[3\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__and4_2
X_10964_ _06905_ _07198_ _07300_ net531 vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12703_ net1989 net263 net383 vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16471_ clknet_leaf_84_wb_clk_i _02225_ _00454_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13683_ team_01_WB.instance_to_wrap.cpu.c0.count\[9\] _04105_ vssd1 vssd1 vccd1 vccd1
+ _04106_ sky130_fd_sc_hd__and2_1
X_10895_ net528 _07234_ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__or2_1
XANTENNA__08692__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15170__A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15422_ net1248 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ net1765 net241 net391 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15353_ net1258 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13402__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12565_ net2225 net204 net399 vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14304_ net1357 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11516_ net1647 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] net877 vssd1 vssd1
+ vccd1 vccd1 _03333_ sky130_fd_sc_hd__mux2_1
X_18072_ net1572 vssd1 vssd1 vccd1 vccd1 la_data_out[114] sky130_fd_sc_hd__buf_2
XFILLER_0_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15284_ net1267 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__inv_2
X_12496_ net3029 net210 net409 vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17023_ clknet_leaf_26_wb_clk_i _02710_ _01006_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14235_ net1367 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11447_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] _07673_ net326 vssd1 vssd1 vccd1
+ vccd1 _07748_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10539__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09608__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14166_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[4\] _04188_ net1695 vssd1
+ vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11200__B2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11378_ _04475_ _07706_ vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__nor2_2
XANTENNA__08512__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ net93 net846 net631 net1919 vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__a22o_1
X_10329_ _06646_ _06653_ _06668_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_52_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[101\] _04254_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[117\]
+ _04383_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_52_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ net1613 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
X_13048_ net1673 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[46\] net853 vssd1 vssd1
+ vccd1 vccd1 _02077_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09046__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1250 net1253 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__buf_4
Xfanout1261 net1269 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__buf_2
X_17856_ clknet_leaf_75_wb_clk_i net1787 _01796_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[126\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1272 net1273 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11476__A1_N net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1283 net1286 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1294 net1303 vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08885__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16807_ clknet_leaf_124_wb_clk_i _02494_ _00790_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09343__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17787_ clknet_leaf_70_wb_clk_i _03463_ _01727_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14999_ net1199 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16738_ clknet_leaf_34_wb_clk_i _02425_ _00721_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08407__A_N _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08132__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16669_ clknet_leaf_49_wb_clk_i _02356_ _00652_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_46_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11812__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09210_ net1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[17\] net936
+ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[14\] net652 _05458_ _05473_
+ _05479_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12767__A1 _07171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17685__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10778__A0 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09072_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[12\] net656 _05385_
+ _05391_ net708 vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_66_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12519__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08023_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] team_01_WB.instance_to_wrap.cpu.f0.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12643__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold700 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold711 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[87\] vssd1 vssd1 vccd1 vccd1
+ net2327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 net2338
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09396__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold733 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[122\] vssd1 vssd1 vccd1 vccd1
+ net2349 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09935__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold744 team_01_WB.instance_to_wrap.cpu.f0.num\[30\] vssd1 vssd1 vccd1 vccd1 net2360
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_64_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold766 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[114\] vssd1 vssd1 vccd1 vccd1
+ net2382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold777 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ net547 net535 net521 net532 vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__o31a_1
Xhold799 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14141__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ _05076_ net558 vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_110_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1400 _03429_ vssd1 vssd1 vccd1 vccd1 net3016 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13495__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1411 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net3027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3038 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15255__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1433 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3049 sky130_fd_sc_hd__dlygate4sd3_1
X_08856_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[3\] net674 net648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1444 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3071 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08795__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09253__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1466 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1477 _02142_ vssd1 vssd1 vccd1 vccd1 net3093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1488 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3104 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout743_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08787_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[0\] net923 vssd1
+ vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1499 team_01_WB.instance_to_wrap.cpu.K0.code\[6\] vssd1 vssd1 vccd1 vccd1 net3115
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13652__C1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09320__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16902__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout910_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09408_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[27\] net689 net657 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[27\]
+ _05747_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10680_ _05901_ _06825_ _06827_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12758__A1 _07111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09339_ net1105 net713 net594 vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09623__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_78_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08316__B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12350_ net2591 net300 net429 vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__mux2_1
XANTENNA__10233__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11430__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11301_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] _05153_ _05154_ vssd1
+ vssd1 vccd1 vccd1 _07641_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_75_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12281_ net1893 net285 net438 vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__mux2_1
XANTENNA__12553__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14020_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[122\] _04250_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[74\]
+ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__a22o_1
X_11232_ _06935_ _07261_ vssd1 vssd1 vccd1 vccd1 _07572_ sky130_fd_sc_hd__nor2_1
XANTENNA__09387__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17408__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08332__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12930__A1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ _07210_ _07255_ net514 vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_36_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10114_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[6\] net820 _04634_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__a22o_1
XANTENNA__14132__B1 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11094_ _07432_ _07433_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__nand2b_1
X_15971_ net1403 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__inv_2
XANTENNA__16432__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17710_ clknet_leaf_102_wb_clk_i _03394_ _01651_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14922_ net1276 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
X_10045_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[0\] net800 net779 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[0\]
+ _06379_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold60 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[15\] vssd1 vssd1 vccd1 vccd1
+ net1676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold71 _03502_ vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17641_ clknet_leaf_114_wb_clk_i _03326_ _01582_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold82 net128 vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
X_14853_ net1209 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__inv_2
Xhold93 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[127\] vssd1 vssd1 vccd1 vccd1
+ net1709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13804_ _04158_ _01834_ _01835_ _01833_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__or4_1
XFILLER_0_118_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17572_ clknet_leaf_61_wb_clk_i _03259_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14784_ net1306 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__inv_2
X_11996_ net2741 net217 net469 vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__mux2_1
XANTENNA__16582__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16523_ clknet_leaf_116_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[21\]
+ _00506_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13735_ _04563_ _04574_ _04503_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__a21oi_1
X_10947_ _06904_ _07281_ _07274_ _07271_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08665__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16454_ clknet_leaf_14_wb_clk_i _02208_ _00437_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13666_ team_01_WB.instance_to_wrap.a1.WRITE_I team_01_WB.instance_to_wrap.a1.READ_I
+ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10878_ _07037_ _07039_ net519 vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15405_ net1207 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12617_ net2373 net305 net398 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__mux2_1
XANTENNA__12749__B2 _03593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16385_ clknet_leaf_65_wb_clk_i _02139_ _00368_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[108\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_22_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13597_ net982 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] _04039_ _04040_
+ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15336_ net1287 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12548_ net2615 net298 net406 vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18055_ net1555 vssd1 vssd1 vccd1 vccd1 la_data_out[97] sky130_fd_sc_hd__buf_2
XFILLER_0_13_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15267_ net1187 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__inv_2
XANTENNA__12463__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ net2027 net285 net414 vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__mux2_1
XANTENNA__14244__A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_2 _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17006_ clknet_leaf_6_wb_clk_i _02693_ _00989_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14218_ net3112 vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09917__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15198_ net1271 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__inv_2
XANTENNA__11185__B1 _07524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12921__A1 _05528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14149_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[55\] _04262_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[23\]
+ _04152_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__a221o_1
Xfanout509 _06032_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14123__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08710_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[5\] net925 vssd1
+ vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__and3_1
XANTENNA__11807__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17908_ net1600 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_0_94_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09690_ _06019_ _06024_ _06029_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__or3_4
XFILLER_0_83_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1080 net1089 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__dlymetal6s2s_1
X_08641_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[10\] net923 vssd1
+ vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__and3_1
Xfanout1091 net1092 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__buf_1
XANTENNA__16925__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17839_ clknet_leaf_63_wb_clk_i _03515_ _01779_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[109\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09504__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15803__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08572_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[19\] net660 _04909_
+ _04910_ _04911_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_136_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08656__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_112_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12638__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10463__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11660__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1066_A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[14\] _04799_
+ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__and3_1
XANTENNA__10215__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09055_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[12\] net898
+ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__and3_1
XANTENNA__12373__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1233_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09369__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08006_ team_01_WB.instance_to_wrap.cpu.f0.state\[2\] vssd1 vssd1 vccd1 vccd1 _04503_
+ sky130_fd_sc_hd__inv_2
Xhold530 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08152__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout693_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold541 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold563 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16455__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold574 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08041__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold585 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[17\] vssd1 vssd1 vccd1 vccd1 net2212
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17700__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14114__B1 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__A team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09957_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[3\] net963 vssd1
+ vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout860_A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[2\] net696 _05225_ _05241_
+ _05242_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__a2111o_1
X_09888_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[5\] net978 vssd1
+ vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__and3_1
Xhold1230 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1241 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 _03481_ vssd1 vssd1 vccd1 vccd1 net2868 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[1\] net688 _05161_ _05167_
+ net708 vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1263 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2879 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1274 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1285 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 net2901
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1296 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2912 sky130_fd_sc_hd__dlygate4sd3_1
X_11850_ net2767 net302 net489 vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ net527 _06972_ _07140_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_16_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11781_ net2458 net283 net497 vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__mux2_1
XANTENNA__12548__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13640__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13520_ _03851_ _03943_ _03850_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__a21oi_1
X_10732_ _05781_ _05898_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__nor2_1
XANTENNA__08327__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13451_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _05381_ _05419_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__a22o_1
X_10663_ _07001_ _07002_ net542 vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__mux2_1
X_12402_ net3085 net272 net422 vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16170_ clknet_leaf_90_wb_clk_i _00012_ _00158_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10594_ net553 _06902_ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__nor2_2
X_13382_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] _05803_ vssd1 vssd1
+ vccd1 vccd1 _03843_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09072__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15121_ net1293 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__inv_2
XANTENNA__08280__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10757__A3 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12333_ net3237 net207 net427 vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12283__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09158__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15052_ net1184 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12264_ net3099 net247 net437 vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__mux2_1
XANTENNA__14999__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14003_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[25\] _04243_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[73\]
+ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__a22o_1
XANTENNA__12903__A1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11706__A2 _07531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08032__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215_ _06750_ _06817_ _06822_ vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10914__A0 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17380__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12195_ net1993 _07838_ net445 vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__mux2_1
XANTENNA__14105__B1 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09780__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _06920_ _07241_ _07275_ _07238_ vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__o211a_1
XANTENNA__16948__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XANTENNA__11627__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13408__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15954_ net1391 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__inv_2
X_11077_ net505 _04919_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__and2b_1
X_10028_ net561 net552 net535 vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__o21ai_1
X_14905_ net1305 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15885_ net1405 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__inv_2
XANTENNA__15623__A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17624_ clknet_leaf_112_wb_clk_i _03309_ _01565_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_14836_ net1287 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__inv_2
XANTENNA__13616__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17555_ clknet_leaf_136_wb_clk_i _03242_ _01538_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14767_ net1215 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__inv_2
XANTENNA__12458__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11979_ net2356 net287 net473 vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__mux2_1
X_16506_ clknet_leaf_109_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[4\]
+ _00489_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13718_ _04105_ net2801 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[8\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_1395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17486_ clknet_leaf_5_wb_clk_i _03173_ _01469_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14698_ net1344 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16437_ clknet_leaf_27_wb_clk_i _02191_ _00420_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13649_ net727 _07507_ net983 vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16368_ clknet_leaf_73_wb_clk_i net1665 _00351_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18107_ net1591 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_125_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15319_ net1199 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12193__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16478__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16299_ clknet_leaf_56_wb_clk_i _02053_ _00282_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08810__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17723__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18038_ net1538 vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__buf_2
XFILLER_0_78_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13552__D1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout306 _07935_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_2
X_09811_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[14\] net773 net738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout317 _07939_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__buf_1
XANTENNA__11173__A3 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout339 _06903_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09742_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[20\] net958
+ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__and3_1
XANTENNA__09523__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09673_ net1120 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[22\] net941
+ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__and3_1
XANTENNA__08877__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08624_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[11\] net677 net662 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[11\]
+ _04954_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__a221o_1
XANTENNA__13607__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09531__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[19\] net655 net653 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[19\]
+ _04894_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12368__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_A _07962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08629__A2 _04968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1183_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13622__A2 _07531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10436__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12830__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08486_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[23\] net934
+ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17253__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12892__A _05678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1350_A net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout706_A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__A team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11397__B1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09107_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[13\] net648 _05428_
+ _05435_ _05437_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_116_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13138__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11301__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09038_ _05264_ _05265_ _05302_ _05377_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_131_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15708__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11020__B net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold360 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[75\] vssd1 vssd1 vccd1 vccd1
+ net1976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[13\] vssd1 vssd1 vccd1 vccd1
+ net1987 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12897__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold382 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _06974_ _06975_ _06883_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_44_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout840 net842 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout851 _03731_ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout862 net863 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_2
Xfanout873 _00017_ vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09514__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout895 _04793_ vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_2
X_12951_ net1803 net873 net360 _03710_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a22o_1
XANTENNA__10124__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08868__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11321__B1 _04534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1060 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2687 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15443__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11902_ net1797 net204 net479 vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1082 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 net2698
+ sky130_fd_sc_hd__dlygate4sd3_1
X_15670_ net1201 vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__inv_2
Xhold1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12882_ net3102 net870 net357 _03662_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__a22o_1
XANTENNA__08983__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14621_ net1365 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__inv_2
X_11833_ net2778 net211 net488 vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__mux2_1
XANTENNA__12278__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13613__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17340_ clknet_leaf_32_wb_clk_i _03027_ _01323_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14552_ net1383 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__inv_2
XANTENNA__10427__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12821__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11764_ net2731 net249 net497 vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13503_ net981 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] _03961_ _03962_
+ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10715_ net553 _06928_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__nand2_1
X_17271_ clknet_leaf_136_wb_clk_i _02958_ _01254_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14483_ net1407 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__inv_2
X_11695_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[12\] net717 vssd1 vssd1 vccd1
+ vccd1 _07893_ sky130_fd_sc_hd__or2_1
XANTENNA__11910__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17746__CLK clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16222_ clknet_leaf_106_wb_clk_i net2037 _00210_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13377__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13434_ _03893_ _03894_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__or2_1
X_10646_ net509 net508 net543 vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11388__B1 _07699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13410__B _05220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16153_ clknet_leaf_98_wb_clk_i _01916_ _00141_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13365_ net585 _07683_ _03834_ net564 _04485_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_51_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10577_ _04741_ _04744_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__or2_2
XFILLER_0_126_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap1168 _07786_ vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__clkbuf_2
X_15104_ net1241 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ net2414 net279 net431 vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16084_ clknet_leaf_102_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[6\]
+ _00072_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16770__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13296_ _07650_ _03779_ _03781_ net825 net1624 vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__o32a_1
XFILLER_0_122_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15035_ net1181 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__inv_2
X_12247_ net3005 net252 net440 vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12178_ net3144 net227 net449 vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__mux2_1
XANTENNA__08520__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11129_ _07466_ _07468_ net553 vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16986_ clknet_leaf_60_wb_clk_i _02673_ _00969_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15937_ net1338 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__inv_2
XANTENNA__09054__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10666__A2 _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15868_ net1345 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__inv_2
XANTENNA__16150__CLK clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08893__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17607_ clknet_leaf_72_wb_clk_i _03294_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_14819_ net1176 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__inv_2
XANTENNA__12188__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15799_ net1354 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__inv_2
X_08340_ net1131 net947 vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__and2_2
XFILLER_0_8_1288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17538_ clknet_leaf_36_wb_clk_i _03225_ _01521_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08271_ net2248 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] net1044 vssd1 vssd1
+ vccd1 vccd1 _03416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17469_ clknet_leaf_49_wb_clk_i _03156_ _01452_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11091__A2 _06882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11820__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10051__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12651__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12879__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09744__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_A _03568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_A _07947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07986_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1 _04484_
+ sky130_fd_sc_hd__inv_2
XANTENNA__14096__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09725_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] net625 _06063_ _06064_
+ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout656_A _04817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1398_A net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] net625 _05994_ _05995_
+ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _04944_ _04945_ _04755_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__mux2_4
XFILLER_0_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12098__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout823_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09587_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[25\] net737 _05908_ _05910_
+ _05914_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_136_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16643__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17769__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08538_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[18\] net691 _04849_ _04863_
+ net706 vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10200__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09275__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08078__A3 _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11015__B net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12826__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08469_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[23\] net897 vssd1
+ vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__and3_1
XANTENNA__11730__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10500_ net1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[31\] net966
+ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__and3b_1
XFILLER_0_68_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09027__A2 _04771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11480_ net367 _07767_ net1983 net874 vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__14020__A2 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16793__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10431_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[27\] net748 net737 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09983__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ net126 net843 net840 net1857 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10362_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[17\] net815 net794 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09139__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10593__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12101_ net1879 net202 net455 vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17149__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13081_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[13\]
+ net854 vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__mux2_1
XANTENNA__12561__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10293_ _06627_ _06628_ _06632_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08978__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ net2402 net211 net465 vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__mux2_1
Xhold190 _02134_ vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13531__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11685__B net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16840_ clknet_leaf_22_wb_clk_i _02527_ _00823_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17299__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout670 net671 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_8
Xfanout681 net682 vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__buf_6
X_16771_ clknet_leaf_20_wb_clk_i _02458_ _00754_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout692 _04772_ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_8
X_13983_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[112\] _04261_ _04262_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[48\]
+ _04274_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__a221o_1
XANTENNA__13295__B1 _04621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15722_ net1273 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11905__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12934_ _05415_ _07757_ _03694_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_18_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09171__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15653_ net1209 vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12865_ net2749 net291 net382 vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
XANTENNA__13405__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09602__C net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14604_ net1330 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__inv_2
XANTENNA__13598__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11816_ net1914 net281 net493 vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__mux2_1
X_15584_ net1241 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__inv_2
XANTENNA__09266__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12796_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] net1056 net364 _03625_
+ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17323_ clknet_leaf_5_wb_clk_i _03010_ _01306_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14535_ net1332 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10805__C1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11747_ net1954 net307 net502 vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__mux2_1
XANTENNA__12270__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17254_ clknet_leaf_40_wb_clk_i _02941_ _01237_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14466_ net1386 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08515__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11678_ _07878_ _07879_ net614 vssd1 vssd1 vccd1 vccd1 _07880_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_133_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14011__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16205_ clknet_leaf_105_wb_clk_i _01965_ _00193_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_133_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13417_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] _05112_ vssd1 vssd1 vccd1
+ vccd1 _03878_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_12_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17185_ clknet_leaf_48_wb_clk_i _02872_ _01168_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10629_ net540 _06968_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_12_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14397_ net1315 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10033__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09974__B1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16136_ clknet_leaf_108_wb_clk_i _00010_ _00124_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13348_ net566 _07680_ _03819_ _03821_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09049__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16067_ clknet_leaf_118_wb_clk_i _01860_ _00055_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12471__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10780__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13279_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] _03753_ vssd1 vssd1 vccd1 vccd1
+ _03768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08888__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15018_ net1279 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__inv_2
XANTENNA__13522__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16516__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11595__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11533__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14078__A2 _04236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16969_ clknet_leaf_10_wb_clk_i _02656_ _00952_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16666__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11815__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[29\] net954
+ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__and3_1
XANTENNA__09081__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09441_ _05779_ _05780_ net598 vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__mux2_2
XFILLER_0_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13589__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09372_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[26\] net657 net656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[26\]
+ _05711_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__a221o_1
XANTENNA__09257__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08323_ net990 net947 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12261__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10955__A _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12646__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08254_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[27\] net3050 net1051 vssd1 vssd1
+ vccd1 vccd1 _03433_ sky130_fd_sc_hd__mux2_1
XANTENNA__14002__A2 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16046__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08185_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[96\] net1686 net1038 vssd1 vssd1
+ vccd1 vccd1 _03502_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout404_A _03565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12381__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1313_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16196__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13513__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08798__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09256__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout773_A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14069__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07969_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 _04467_
+ sky130_fd_sc_hd__inv_2
XANTENNA__11725__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09708_ net1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[21\] net941
+ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__and3_1
X_10980_ net531 _07182_ _07319_ net376 vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__a22o_1
XANTENNA__10849__B _06472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09639_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[23\] net948
+ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_84_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08319__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11026__A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12650_ net2858 net307 net393 vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09248__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11601_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\]
+ _07817_ vssd1 vssd1 vccd1 vccd1 _07818_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12581_ net2665 net298 net402 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12556__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ net1356 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11532_ net1890 net1157 net587 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[21\] vssd1
+ vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08335__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14056__B _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_830 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire323 _07352_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12004__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ net1354 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13201__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11463_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[15\] _07755_ _07758_ vssd1 vssd1
+ vccd1 vccd1 _07759_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10015__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13202_ net6 net836 net628 net1721 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__o22a_1
X_10414_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[27\] net970
+ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__and3_1
X_14182_ net1807 _04452_ net1169 vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11394_ net1062 _07668_ _07714_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1
+ vssd1 vccd1 vccd1 _07720_ sky130_fd_sc_hd__a31o_1
X_13133_ net76 net848 net632 net3209 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10345_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[17\] net953
+ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09166__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13064_ net1625 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[30\] net858 vssd1 vssd1
+ vccd1 vccd1 _02061_ sky130_fd_sc_hd__mux2_1
X_17941_ net1441 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XANTENNA__10318__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10276_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[19\] net746 _06613_ _06614_
+ _06615_ vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1410 net1413 vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__buf_2
X_12015_ net2670 net283 net469 vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__mux2_1
X_17872_ clknet_leaf_91_wb_clk_i _03547_ _01812_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16823_ clknet_leaf_140_wb_clk_i _02510_ _00806_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13966_ _04238_ _04257_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__nor2_8
X_16754_ clknet_leaf_134_wb_clk_i _02441_ _00737_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15705_ net1259 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__inv_2
X_12917_ _05564_ net577 vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16685_ clknet_leaf_140_wb_clk_i _02372_ _00668_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13897_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\] _04141_ vssd1 vssd1 vccd1
+ vccd1 _04200_ sky130_fd_sc_hd__or2_1
XANTENNA__11061__A1_N _05042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15636_ net1288 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12848_ net2277 net268 net380 vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__mux2_1
XANTENNA__09239__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16069__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15567_ net1217 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__inv_2
XANTENNA__12466__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12779_ net1762 net641 net608 _03614_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a22o_1
XANTENNA__17314__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08998__A1 _05337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17306_ clknet_leaf_59_wb_clk_i _02993_ _01289_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14518_ net1335 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15498_ net1282 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17237_ clknet_leaf_124_wb_clk_i _02924_ _01220_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14449_ net1378 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold904 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
X_17168_ clknet_leaf_13_wb_clk_i _02855_ _01151_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold915 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[112\] vssd1 vssd1 vccd1 vccd1
+ net2531 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09411__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold926 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[104\] vssd1 vssd1 vccd1 vccd1
+ net2542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16119_ clknet_leaf_109_wb_clk_i _01894_ _00107_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold937 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[32\] vssd1 vssd1 vccd1 vccd1
+ net2564 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09990_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[2\] net805 net751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold959 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[111\] vssd1 vssd1 vccd1 vccd1
+ net2575 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17099_ clknet_leaf_144_wb_clk_i _02786_ _01082_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08941_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[6\] net917 vssd1
+ vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09507__C net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09175__A1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[3\] net664 _05198_ _05200_
+ _05202_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__a2111o_1
Xhold1604 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1615 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1626 _03449_ vssd1 vssd1 vccd1 vccd1 net3242 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1637 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3253 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3264 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1659 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3275 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout187_A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09478__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout354_A _03741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1096_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09424_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[28\] net689 net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[28\]
+ _05763_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_118_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09355_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[25\] net670 net651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__a22o_1
XANTENNA__12376__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10685__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10245__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08306_ net1132 net965 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__and2_2
XANTENNA_clkbuf_leaf_68_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_118_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12785__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09286_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[22\] net886 vssd1
+ vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17807__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08237_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[44\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[36\]
+ net1041 vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07994__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08168_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[113\] net1680 net1052 vssd1 vssd1
+ vccd1 vccd1 _03519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10548__A1 _06098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09402__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout890_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_108_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout988_A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08610__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08099_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[0\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10130_ _06438_ _06440_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__nor2_1
X_10061_ _06369_ _06400_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_86_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13820_ net1721 net833 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[13\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_86_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13751_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _04140_
+ sky130_fd_sc_hd__nand3_1
X_10963_ net542 _06940_ _06942_ _07302_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_67_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16211__CLK clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13670__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12702_ net2529 net268 net383 vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__mux2_1
X_16470_ clknet_leaf_84_wb_clk_i _02224_ _00453_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13682_ team_01_WB.instance_to_wrap.cpu.c0.count\[8\] team_01_WB.instance_to_wrap.cpu.c0.count\[7\]
+ _04103_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10894_ _07137_ _07181_ net514 vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15421_ net1262 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__inv_2
X_12633_ net3201 net272 net393 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__mux2_1
XANTENNA__12286__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14067__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10595__A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10236__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15352_ net1178 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__inv_2
XANTENNA__11433__C1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12564_ net2053 net206 net399 vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17487__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09641__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14303_ net1353 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11515_ net2019 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] net877 vssd1 vssd1
+ vccd1 vccd1 _03334_ sky130_fd_sc_hd__mux2_1
X_18071_ net1571 vssd1 vssd1 vccd1 vccd1 la_data_out[113] sky130_fd_sc_hd__buf_2
X_15283_ net1281 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12495_ net3171 net250 net409 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17022_ clknet_leaf_44_wb_clk_i _02709_ _01005_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09929__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14234_ net1364 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__inv_2
X_11446_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] _07674_ _07747_ vssd1 vssd1 vccd1
+ vccd1 _03367_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14165_ _04195_ _04443_ net1412 vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08601__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11377_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] _07705_ vssd1 vssd1 vccd1 vccd1
+ _07706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13116_ net1916 net843 net631 team_01_WB.instance_to_wrap.a1.ADR_I\[27\] vssd1 vssd1
+ vccd1 vccd1 _02025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10328_ _06657_ _06659_ _06663_ _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__or4_1
X_14096_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[69\] _04233_ _04253_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ net1612 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_124_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ net2345 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[47\] net861 vssd1 vssd1
+ vccd1 vccd1 _02078_ sky130_fd_sc_hd__mux2_1
X_10259_ _06193_ _06218_ _06192_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1240 net1245 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1251 net1253 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__buf_4
X_17855_ clknet_leaf_63_wb_clk_i _03531_ _01795_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[125\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout1262 net1265 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__buf_4
Xfanout1273 net1303 vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__clkbuf_4
Xfanout1284 net1286 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__buf_4
X_16806_ clknet_leaf_42_wb_clk_i _02493_ _00789_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1295 net1302 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17786_ clknet_leaf_76_wb_clk_i _03462_ _01726_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_14998_ net1247 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__inv_2
XANTENNA_wire322_A _07464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16737_ clknet_leaf_41_wb_clk_i _02424_ _00720_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09062__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13949_ _04218_ _04229_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__nor2_4
XFILLER_0_18_1344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_102_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16668_ clknet_leaf_32_wb_clk_i _02355_ _00651_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15619_ net1177 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__inv_2
XANTENNA__12196__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16599_ clknet_leaf_118_wb_clk_i _02286_ _00582_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09140_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[14\] net699 _05461_
+ _05462_ _05468_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_57_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09071_ _05407_ _05408_ _05409_ _05410_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16854__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08022_ _04505_ _04516_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__or2_2
XFILLER_0_115_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold701 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[106\] vssd1 vssd1 vccd1 vccd1
+ net2328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11727__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold723 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09396__A1 _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13192__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold734 _03528_ vssd1 vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold745 team_01_WB.instance_to_wrap.a1.ADR_I\[31\] vssd1 vssd1 vccd1 vccd1 net2361
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold767 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[91\] vssd1 vssd1 vccd1 vccd1
+ net2383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold778 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[54\] vssd1 vssd1 vccd1 vccd1
+ net2394 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] net627 _06311_ _06312_
+ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__a22o_4
XFILLER_0_42_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold789 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10950__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08924_ net547 net535 net532 net521 vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__or4_4
XFILLER_0_42_1673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1011_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_141_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1401 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3017 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09534__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[3\] net916 vssd1
+ vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__and3_1
Xhold1412 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1423 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 net3039
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout471_A _07952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1434 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[19\] vssd1 vssd1 vccd1 vccd1
+ net3050 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16234__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1445 team_01_WB.instance_to_wrap.cpu.DM0.state\[0\] vssd1 vssd1 vccd1 vccd1 net3061
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout569_A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1456 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3072 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08786_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[0\] net885 vssd1
+ vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__and3_1
Xhold1467 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1478 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net3094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1489 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3105 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12455__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout736_A _04687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1380_A net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09320__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15271__A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07989__A team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09871__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09407_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[27\] net661 net656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09700__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout903_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09338_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] net704 _05672_ _05677_
+ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__o22a_4
XANTENNA__10769__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09269_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[20\] net673 net656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[20\]
+ _05608_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12834__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11300_ _05153_ _05154_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1
+ vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_75_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12280_ net2638 net251 net436 vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__mux2_1
XANTENNA__11958__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09387__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11231_ _07569_ _07570_ vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08332__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11162_ _07382_ _07501_ _07042_ _07101_ vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_120_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10113_ _06449_ _06450_ _06451_ _06452_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_8_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15970_ net1391 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__inv_2
X_11093_ net535 _06366_ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08986__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09444__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14921_ net1215 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
X_10044_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[0\] net753 _06373_ _06383_
+ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_69_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12694__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold50 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[9\] vssd1 vssd1 vccd1 vccd1
+ net1666 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold61 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[10\] vssd1 vssd1 vccd1 vccd1
+ net1688 sky130_fd_sc_hd__dlygate4sd3_1
X_17640_ clknet_leaf_113_wb_clk_i _03325_ _01581_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_14852_ net1237 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__inv_2
Xhold83 _01994_ vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 _03533_ vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16727__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13803_ _04159_ _04181_ _04182_ _04154_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a22o_1
X_17571_ clknet_leaf_61_wb_clk_i _03258_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14783_ net1306 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__inv_2
X_11995_ net2067 net221 net469 vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11913__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10457__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16522_ clknet_leaf_116_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[20\]
+ _00505_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13734_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] _04516_ _04524_ _04134_ vssd1
+ vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10946_ _07284_ _07285_ net519 vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09862__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13665_ net982 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] _04095_ _04096_
+ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a22o_1
X_16453_ clknet_leaf_23_wb_clk_i _02207_ _00436_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10877_ net555 _07216_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16877__CLK clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10209__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11214__A _07171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12616_ net2226 net311 net396 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__mux2_1
XANTENNA__12749__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15404_ net1181 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__inv_2
X_16384_ clknet_leaf_73_wb_clk_i net2497 _00367_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13596_ net723 _07188_ net1068 vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__o21a_1
XANTENNA__09614__A2 _04636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15335_ net1300 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12547_ net2153 net280 net404 vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18054_ net1554 vssd1 vssd1 vccd1 vccd1 la_data_out[96] sky130_fd_sc_hd__buf_2
XFILLER_0_123_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15266_ net1266 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__inv_2
X_12478_ net3224 net251 net412 vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__mux2_1
XANTENNA_3 _05490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08523__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13174__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17005_ clknet_leaf_140_wb_clk_i _02692_ _00988_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14217_ net3034 vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11429_ net326 _07738_ _07739_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_1624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15197_ net1253 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11185__B2 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10491__C net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14148_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[15\] _04226_ _04260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[63\]
+ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09057__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17502__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14079_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[28\] _04243_ _04245_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[84\]
+ _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17907_ net1599 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XANTENNA__08896__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12685__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1070 net1071 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__buf_2
X_08640_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[10\] net888
+ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__and3_1
Xfanout1081 net1082 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_2
X_17838_ clknet_leaf_64_wb_clk_i _03514_ _01778_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[108\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout1092 net1095 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__buf_2
XFILLER_0_94_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08571_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[19\] net900 vssd1
+ vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__and3_1
X_17769_ clknet_leaf_78_wb_clk_i _03445_ _01709_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13634__B1 team_01_WB.instance_to_wrap.cpu.IM0.pc_enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11823__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15091__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08417__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09123_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[14\] net925
+ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout317_A _07939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1059_A team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09054_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[12\] net895 vssd1
+ vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09529__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17032__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08433__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08005_ team_01_WB.instance_to_wrap.cpu.c0.count\[16\] vssd1 vssd1 vccd1 vccd1 _04502_
+ sky130_fd_sc_hd__inv_2
Xhold520 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1226_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold542 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold553 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08041__A1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold564 team_01_WB.instance_to_wrap.a1.ADR_I\[4\] vssd1 vssd1 vccd1 vccd1 net2180
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold575 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold586 team_01_WB.instance_to_wrap.cpu.f0.num\[10\] vssd1 vssd1 vccd1 vccd1 net2202
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A _04780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold597 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17182__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08592__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[3\] net960 vssd1
+ vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__and3_1
XANTENNA__08579__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08907_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[2\] net880 vssd1
+ vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09887_ net993 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[5\] net963 vssd1
+ vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout853_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1220 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1231 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2847 sky130_fd_sc_hd__dlygate4sd3_1
X_08838_ _05175_ _05176_ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__or3_1
Xhold1242 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2858 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10203__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1253 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[27\] vssd1 vssd1 vccd1 vccd1
+ net2869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2880 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10151__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1275 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1286 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2902 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11018__B _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ _05105_ _05106_ _05107_ _05108_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__or4_1
Xhold1297 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10800_ net523 _07139_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__nand2_1
XANTENNA__10439__B1 _06777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ net2473 net251 net496 vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_3__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09844__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08608__A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10731_ _05115_ _07069_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08327__B net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11034__A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13450_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _04946_ _03910_ vssd1
+ vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__o21a_1
X_10662_ _06526_ net340 net546 vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14050__B1 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12401_ net3164 net243 net419 vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_123_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12564__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] _05803_ vssd1 vssd1
+ vccd1 vccd1 _03842_ sky130_fd_sc_hd__or2_1
X_10593_ net555 _06930_ _06931_ _06932_ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_23_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15120_ net1270 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__inv_2
X_12332_ net2657 net275 net429 vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08343__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15051_ net1297 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12263_ net3152 net213 net437 vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14002_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[49\] _04262_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11214_ _07171_ _07207_ _07251_ _07542_ vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08032__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12194_ net3234 net218 net445 vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__mux2_1
XANTENNA__10914__A1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11908__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11145_ _05263_ _07484_ vssd1 vssd1 vccd1 vccd1 _07485_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
X_15953_ net1333 vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__inv_2
XANTENNA__13408__B _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17675__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ _04884_ _06672_ _07127_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09605__C net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ net561 net552 net534 vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__or3_1
XANTENNA__11209__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10678__B1 _07016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14904_ net1171 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
X_15884_ net1386 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__inv_2
XANTENNA__10142__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17623_ clknet_leaf_111_wb_clk_i _03308_ _01564_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_14835_ net1280 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11643__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13424__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17554_ clknet_leaf_129_wb_clk_i _03241_ _01537_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14766_ net1284 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__inv_2
X_11978_ net2258 net256 net472 vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__mux2_1
XANTENNA__13092__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09835__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08518__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16505_ clknet_leaf_108_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[3\]
+ _00488_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10929_ net563 _07253_ _07264_ _07268_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__a211o_2
X_13717_ team_01_WB.instance_to_wrap.cpu.c0.count\[7\] _04103_ net2800 vssd1 vssd1
+ vccd1 vccd1 _04128_ sky130_fd_sc_hd__a21oi_1
X_14697_ net1343 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__inv_2
X_17485_ clknet_leaf_140_wb_clk_i _03172_ _01468_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16436_ clknet_leaf_104_wb_clk_i _02190_ _00419_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13648_ net188 _04081_ _04082_ net727 vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__a211o_1
XFILLER_0_27_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16367_ clknet_leaf_67_wb_clk_i _02121_ _00350_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12474__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13579_ _03917_ _04024_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14255__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18106_ net636 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08271__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15318_ net1198 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__inv_2
X_16298_ clknet_leaf_61_wb_clk_i _02052_ _00281_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[21\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_124_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18037_ net1537 vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__buf_2
XFILLER_0_83_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15249_ net1292 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09810_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[14\] net815 net749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__a22o_1
XANTENNA__11818__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout307 _07935_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_2
XANTENNA__11169__C_N _07308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__B2 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout318 net321 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_2
Xfanout329 _07101_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10381__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13304__C1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09084__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[20\] net952
+ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__and3_1
XANTENNA__13318__B net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09672_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[22\] net951
+ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__and3_1
X_08623_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[11\] net684 _04962_
+ net707 vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12649__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout267_A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08554_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[19\] net900
+ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08485_ net1087 net935 vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__and2_2
XFILLER_0_76_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08495__D1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11633__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10841__A0 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1176_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14032__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12384__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout601_A _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16422__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09106_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[13\] net669 _05427_ _05438_
+ _05441_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_131_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09037_ _05006_ _05338_ _05374_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__and3_1
XANTENNA__13138__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11301__B _05153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold350 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold361 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17698__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold372 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14099__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout830 _04578_ vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__buf_2
Xfanout841 net842 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__buf_4
Xfanout852 net853 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__clkbuf_4
X_09939_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] net766 net623 vssd1
+ vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__o21a_1
XANTENNA__12649__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout863 net869 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__buf_2
Xfanout874 net875 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_2
Xfanout885 net886 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__buf_4
XANTENNA__15724__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout896 net897 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__buf_4
X_12950_ net1036 net583 _03709_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10124__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1050 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11321__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold1061 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2677 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11901_ net3044 net207 net479 vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__mux2_1
Xhold1072 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[102\] vssd1 vssd1 vccd1 vccd1
+ net2688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12881_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[28\] _03661_ net1030 vssd1
+ vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__mux2_1
Xhold1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2699 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12559__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14620_ net1360 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__inv_2
X_11832_ net3254 net250 net488 vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__mux2_1
XANTENNA__17078__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08338__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13613__A3 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14551_ net1338 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09160__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11763_ net3227 net213 net497 vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12821__B2 _03643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10714_ net553 _06928_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__and2_2
X_13502_ net724 _07019_ net1067 vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14482_ net1387 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__inv_2
X_17270_ clknet_leaf_1_wb_clk_i _02957_ _01253_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11694_ net2852 net258 net501 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__mux2_1
XANTENNA__14023__B1 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13377__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16221_ clknet_leaf_105_wb_clk_i net1724 _00209_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
X_13433_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] net595 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__a21oi_1
X_10645_ _06098_ net505 net543 vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12294__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16152_ clknet_leaf_97_wb_clk_i _01915_ _00140_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13364_ net1064 net1065 vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__or2_1
X_10576_ net503 _06882_ net370 vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__o21a_1
XANTENNA__09450__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12315_ net2719 _07912_ net432 vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__mux2_1
X_15103_ net1256 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__inv_2
XANTENNA__13129__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16083_ clknet_leaf_102_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[5\]
+ _00071_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13295_ _03751_ _03780_ _04621_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__a21oi_1
X_15034_ net1191 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__inv_2
XANTENNA__13534__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12246_ net2761 net230 net440 vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_91_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12177_ net2379 net290 net450 vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__mux2_1
XANTENNA__10542__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10363__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ net525 _07256_ _07467_ _06906_ vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_78_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16985_ clknet_leaf_58_wb_clk_i _02672_ _00968_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_15936_ net1336 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__inv_2
X_11059_ net557 _06281_ _07384_ _06251_ _05076_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__a32o_1
XANTENNA__10115__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09632__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15867_ net1350 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__inv_2
XANTENNA__12469__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17606_ clknet_leaf_72_wb_clk_i _03293_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14818_ net1266 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__inv_2
XANTENNA__09269__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15798_ net1381 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17537_ clknet_leaf_42_wb_clk_i _03224_ _01520_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12812__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14749_ net1309 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08270_ net2758 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] net1051 vssd1 vssd1
+ vccd1 vccd1 _03417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17468_ clknet_leaf_37_wb_clk_i _03155_ _01451_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16419_ clknet_leaf_86_wb_clk_i _02173_ _00402_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17399_ clknet_leaf_136_wb_clk_i _03086_ _01382_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11402__A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09441__A0 _05779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16595__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08711__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10354__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07985_ team_01_WB.instance_to_wrap.cpu.f0.i\[10\] vssd1 vssd1 vccd1 vccd1 _04483_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout384_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\] net764 net621 vssd1
+ vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10106__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09542__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] net764 net621 vssd1
+ vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__o21a_1
XANTENNA__12379__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout551_A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1293_A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout649_A _04823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08606_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] net619 net593 vssd1 vssd1
+ vccd1 vccd1 _04946_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_2_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[25\] net786 net762 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__a22o_1
XANTENNA__11067__B1 _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08537_ _04873_ _04874_ _04875_ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__nor4_1
XFILLER_0_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12803__B2 _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout816_A _04636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08468_ net1004 net896 vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__and2_4
XANTENNA__14005__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08399_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] net712 net620 _04724_ vssd1
+ vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_45_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11312__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10430_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[27\] net813 _06757_ _06760_
+ _06761_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_33_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09432__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08324__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10361_ _06683_ _06698_ _06699_ _06700_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__or4_1
XFILLER_0_131_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12842__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12100_ net2771 net207 net455 vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__mux2_1
XANTENNA__13516__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13080_ net1717 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[14\] net853 vssd1 vssd1
+ vccd1 vccd1 _02045_ sky130_fd_sc_hd__mux2_1
X_10292_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[19\] net735 _06629_ _06630_
+ _06631_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_108_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12031_ net2647 net248 net465 vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__mux2_1
XANTENNA__08538__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 _02007_ vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1
+ net1807 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08340__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16318__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11542__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout660 _04813_ vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_8
Xfanout671 _04800_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_8
XPHY_EDGE_ROW_69_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16770_ clknet_leaf_34_wb_clk_i _02457_ _00753_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout682 _04787_ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__buf_6
X_13982_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[104\] _04252_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[72\]
+ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__a22o_1
Xfanout693 net694 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08994__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15721_ net1222 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12933_ net359 _03697_ _03698_ net872 net2131 vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a32o_1
X_17969__1469 vssd1 vssd1 vccd1 vccd1 _17969__1469/HI net1469 sky130_fd_sc_hd__conb_1
XANTENNA__12289__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15652_ net1191 vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12864_ net2196 net314 net381 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14603_ net1401 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11815_ net2014 net304 net493 vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15583_ net1254 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__inv_2
X_12795_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[11\] _07207_ net1028 vssd1 vssd1
+ vccd1 vccd1 _03625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11921__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17322_ clknet_leaf_10_wb_clk_i _03009_ _01305_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14534_ net1335 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11746_ _07932_ _07933_ _07934_ net612 vssd1 vssd1 vccd1 vccd1 _07935_ sky130_fd_sc_hd__a22o_2
XFILLER_0_12_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17253_ clknet_leaf_40_wb_clk_i _02940_ _01236_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14465_ net1316 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11677_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] _07811_ vssd1 vssd1
+ vccd1 vccd1 _07879_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_133_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16204_ clknet_leaf_62_wb_clk_i _01964_ _00192_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13416_ _03871_ _03876_ _03870_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__a21o_1
X_10628_ _04706_ _06857_ net545 vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17184_ clknet_leaf_33_wb_clk_i _02871_ _01167_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14396_ net1316 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09423__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09974__A1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16135_ clknet_leaf_107_wb_clk_i _00009_ _00123_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11230__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13347_ net585 _07687_ _03820_ net830 vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10559_ net540 _06896_ _06898_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13507__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16066_ clknet_leaf_118_wb_clk_i _01859_ _00054_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_13278_ _03748_ _03766_ _04518_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09726__A1 _05570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15017_ net1216 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__inv_2
XANTENNA__13522__A2 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ net2992 net219 net441 vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__mux2_1
XANTENNA__11595__C team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11533__B2 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17243__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16968_ clknet_leaf_22_wb_clk_i _02655_ _00951_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10004__C net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15919_ net1410 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__inv_2
XANTENNA__11297__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12199__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16899_ clknet_leaf_18_wb_clk_i _02586_ _00882_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17393__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] net712 _04841_ vssd1 vssd1
+ vccd1 vccd1 _05780_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09371_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[26\] net695 net692 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__a22o_1
XANTENNA__08409__C _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13589__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11831__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_96_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12797__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ net1148 net1151 net1153 net1147 vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__and4b_1
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08706__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10955__B _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08253_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[28\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[20\]
+ net1041 vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13746__C1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08184_ net2423 net2987 net1052 vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13210__A1 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08768__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12662__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1041_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1139_A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09537__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout599_A _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13513__A2 _07088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10327__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11524__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1306_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout766_A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16610__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17736__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1 _04466_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09707_ net1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[21\] net943
+ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__and3_1
XANTENNA__09703__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11307__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09638_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[23\] net951 vssd1
+ vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11026__B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09569_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[25\] net973
+ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12837__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\]
+ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _07814_ vssd1 vssd1 vccd1 vccd1
+ _07817_ sky130_fd_sc_hd__and4_1
X_12580_ net1937 net280 net399 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11531_ net1679 net1157 net587 net1111 vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__a22o_1
XANTENNA__11460__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08335__B net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire324 _07258_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_1
XANTENNA__14056__C _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14250_ net1354 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11462_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] _07757_ net877 vssd1 vssd1
+ vccd1 vccd1 _07758_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_123_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09405__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13201__A1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13201_ net7 net837 net630 net2343 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__a22o_1
X_10413_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[27\] net968
+ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__and3_1
X_14181_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[11\] _04452_ vssd1 vssd1 vccd1
+ vccd1 _04453_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11393_ _04466_ _07715_ _07719_ net325 vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__o211a_1
XANTENNA__12572__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12960__A0 team_01_WB.instance_to_wrap.cpu.f0.write_data\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13132_ net77 net848 net631 net1792 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08989__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17266__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input62_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[17\] net978
+ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13063_ net3182 net2982 net861 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__mux2_1
X_17940_ net1440 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_29_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10275_ net987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[19\] net948 vssd1
+ vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__and3_1
XANTENNA__11515__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12014_ net2295 net254 net467 vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__mux2_1
Xfanout1400 net1401 vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__buf_4
Xfanout1411 net1412 vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__buf_4
X_17871_ clknet_leaf_82_wb_clk_i _03546_ _01811_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16290__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11916__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16822_ clknet_leaf_1_wb_clk_i _02509_ _00805_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout490 _07947_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16753_ clknet_leaf_17_wb_clk_i _02440_ _00736_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13965_ _04219_ _04231_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_31_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15704_ net1178 vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__inv_2
X_12916_ net358 _03685_ _03686_ net871 net2065 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__a32o_1
X_16684_ clknet_leaf_133_wb_clk_i _02371_ _00667_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13896_ _04141_ net571 _04199_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__and3b_1
X_15635_ net1280 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12847_ net2442 net236 net379 vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11651__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13432__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ net1285 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__inv_2
XANTENNA__09644__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08526__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12778_ net365 _03612_ _03613_ net1056 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\]
+ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_44_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ clknet_leaf_55_wb_clk_i _02992_ _01288_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14517_ net1405 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11451__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11729_ net612 _07799_ _07920_ _07919_ vssd1 vssd1 vccd1 vccd1 _07921_ sky130_fd_sc_hd__a31o_2
X_15497_ net1217 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__inv_2
XANTENNA__10494__C net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17236_ clknet_leaf_12_wb_clk_i _02923_ _01219_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14448_ net1376 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12482__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17167_ clknet_leaf_144_wb_clk_i _02854_ _01150_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14379_ net1319 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold905 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14263__A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold916 _03518_ vssd1 vssd1 vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold927 _03510_ vssd1 vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12951__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08899__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16118_ clknet_leaf_100_wb_clk_i _01893_ _00106_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold938 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold949 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
X_17098_ clknet_leaf_2_wb_clk_i _02785_ _01081_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08940_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[6\] net924 vssd1
+ vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__and3_1
XANTENNA__16633__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16049_ clknet_leaf_87_wb_clk_i _01842_ _00037_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_86_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08871_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[3\] _04800_ net652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[3\]
+ _05196_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_131_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1605 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[38\] vssd1 vssd1 vccd1 vccd1
+ net3221 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15094__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1616 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1627 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net3243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1638 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3265 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09092__A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16783__CLK clknet_leaf_143_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18039__1539 vssd1 vssd1 vccd1 vccd1 _18039__1539/HI net1539 sky130_fd_sc_hd__conb_1
X_09423_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[28\] net683 net680 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12657__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout347_A net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1089_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[25\] net701 net650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08436__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08305_ net1146 net1151 net1153 net1149 vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_63_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13982__A2 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[22\] net886
+ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout514_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1256_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[45\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[37\]
+ net1040 vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13195__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08167_ net2382 net2328 net1042 vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12392__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13734__A2 _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17968__1468 vssd1 vssd1 vccd1 vccd1 _17968__1468/HI net1468 sky130_fd_sc_hd__conb_1
XFILLER_0_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12942__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08098_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[4\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[7\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[6\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__or4b_1
XFILLER_0_31_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout883_A _04803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13498__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10060_ _06367_ _06368_ _06366_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11736__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13750_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__nand2_1
X_10962_ net542 _07301_ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09874__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12701_ net2157 net236 net383 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11681__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12567__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13681_ team_01_WB.instance_to_wrap.cpu.c0.count\[7\] _04103_ vssd1 vssd1 vccd1 vccd1
+ _04104_ sky130_fd_sc_hd__nand2_1
X_10893_ _06677_ _07113_ net344 vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15420_ net1173 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12632_ net3181 net243 net391 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__mux2_1
XANTENNA__10595__B _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08346__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16506__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15351_ net1189 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__inv_2
X_12563_ net1885 net277 net401 vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09876__S net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14302_ net1356 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__inv_2
X_11514_ net1639 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] net877 vssd1 vssd1
+ vccd1 vccd1 _03335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18070_ net1570 vssd1 vssd1 vccd1 vccd1 la_data_out[112] sky130_fd_sc_hd__buf_2
X_15282_ net1233 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12494_ net2898 net214 net409 vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17021_ clknet_leaf_21_wb_clk_i _02708_ _01004_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13186__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14233_ net1360 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__inv_2
X_11445_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] _07674_ net326 vssd1 vssd1 vccd1
+ vccd1 _07747_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10539__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11197__C1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12933__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[4\] _04188_ vssd1 vssd1 vccd1
+ vccd1 _04443_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11376_ _04477_ _07704_ vssd1 vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__nor2_1
XANTENNA__09608__C net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08512__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ net1719 net843 net631 team_01_WB.instance_to_wrap.a1.ADR_I\[28\] vssd1 vssd1
+ vccd1 vccd1 _02026_ sky130_fd_sc_hd__a22o_1
X_10327_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[18\] net794 _06664_ _06665_
+ _06666_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_128_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14095_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[29\] _04243_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[109\]
+ _04381_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__a221o_1
XANTENNA__15907__A net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ net1611 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
X_13046_ net2376 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[48\] net868 vssd1 vssd1
+ vccd1 vccd1 _02079_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10258_ _06221_ _06469_ _06472_ _06597_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__or4_4
XFILLER_0_56_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1230 net1231 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__buf_2
XFILLER_0_98_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11646__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1241 net1245 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__buf_4
XANTENNA__13427__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17854_ clknet_leaf_65_wb_clk_i _03530_ _01794_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[124\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__10172__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10189_ _04750_ _05376_ _05006_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1252 net1253 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1263 net1265 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__buf_4
Xfanout1274 net1277 vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__buf_4
Xfanout1285 net1286 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__buf_2
X_16805_ clknet_leaf_37_wb_clk_i _02492_ _00788_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1296 net1302 vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__buf_2
X_17785_ clknet_leaf_77_wb_clk_i net2004 _01725_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09343__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14997_ net1225 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16736_ clknet_leaf_30_wb_clk_i _02423_ _00719_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13948_ _04227_ _04237_ _04239_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__and3_4
XFILLER_0_117_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09865__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09640__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16667_ clknet_leaf_50_wb_clk_i _02354_ _00650_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12477__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11672__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13879_ team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] _03575_ _04136_ _00005_ vssd1
+ vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_read_i sky130_fd_sc_hd__a31o_1
XANTENNA__14258__A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15618_ net1266 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13413__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16186__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16598_ clknet_leaf_117_wb_clk_i _02285_ _00581_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17431__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15549_ net1250 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09070_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[12\] net662 _05387_
+ _05399_ _05402_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_86_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08021_ _04505_ _04516_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17219_ clknet_leaf_19_wb_clk_i _02906_ _01202_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10725__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11727__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold702 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11410__A team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09087__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold713 _03512_ vssd1 vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold724 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold735 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[91\] vssd1 vssd1 vccd1 vccd1
+ net2351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold746 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold757 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 _02130_ vssd1 vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold779 _03468_ vssd1 vssd1 vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09972_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\] net766 net623 vssd1
+ vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__o21a_1
XANTENNA__09148__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ net525 net516 vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__nand2_4
XANTENNA__14141__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08356__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout297_A _07926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1402 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3018 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08854_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[3\] net903 vssd1
+ vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__and3_1
Xhold1413 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3029 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10163__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1004_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1424 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3040 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1435 _03433_ vssd1 vssd1 vccd1 vccd1 net3051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1446 _00013_ vssd1 vssd1 vccd1 vccd1 net3062 sky130_fd_sc_hd__dlygate4sd3_1
X_08785_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[0\] net906 vssd1
+ vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__and3_1
Xhold1457 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net3073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net3084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout464_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1479 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 net3095
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09856__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13652__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16529__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12387__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout631_A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1373_A net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09406_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[27\] net688 _04797_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\]
+ _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09337_ _05661_ _05674_ _05675_ _05676_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16679__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09268_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[20\] net904
+ net657 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[20\] vssd1 vssd1 vccd1
+ vccd1 _05608_ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11430__A3 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13168__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08219_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[62\] net2394 net1042 vssd1 vssd1
+ vccd1 vccd1 _03468_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09199_ net1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[17\] net897
+ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11230_ _05934_ _05965_ _07568_ net344 vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11161_ _05076_ net333 _07500_ net371 vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_82_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12850__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10112_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[6\] net754 net751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__a22o_1
XANTENNA__14132__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11092_ net535 _06366_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_8_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13852__A_N net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14920_ net1276 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
X_10043_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[0\] net817 net791 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold40 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[29\] vssd1 vssd1 vccd1 vccd1
+ net1656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[34\] vssd1 vssd1 vccd1 vccd1 net1667
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[19\] vssd1 vssd1 vccd1 vccd1
+ net1678 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ net1186 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__inv_2
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 team_01_WB.instance_to_wrap.cpu.f0.write_data\[13\] vssd1 vssd1 vccd1 vccd1
+ net1689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[27\] vssd1 vssd1 vccd1 vccd1
+ net1700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[31\] vssd1 vssd1 vccd1 vccd1
+ net1711 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ _01836_ _04164_ _04173_ _01837_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__a31o_1
X_17570_ clknet_leaf_61_wb_clk_i _03257_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09847__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14782_ net1312 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__inv_2
XANTENNA__13643__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11994_ net3070 net226 net467 vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__mux2_1
X_16521_ clknet_leaf_115_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[19\]
+ _00504_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17454__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09311__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13733_ team_01_WB.instance_to_wrap.cpu.DM0.dhit team_01_WB.instance_to_wrap.cpu.f0.state\[3\]
+ team_01_WB.instance_to_wrap.cpu.f0.state\[0\] team_01_WB.EN_VAL_REG vssd1 vssd1
+ vccd1 vccd1 _04134_ sky130_fd_sc_hd__a22o_1
X_10945_ net375 _06158_ net374 net342 net551 net539 vssd1 vssd1 vccd1 vccd1 _07285_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12297__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16452_ clknet_leaf_123_wb_clk_i _02206_ _00435_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13664_ net723 _07489_ net1068 vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10876_ net524 _07215_ _07213_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_112_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15403_ net1297 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12615_ net2642 net294 net398 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__mux2_1
XANTENNA__11214__B _07207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16383_ clknet_leaf_67_wb_clk_i net2600 _00366_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13595_ net187 _04037_ _04038_ net728 vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11957__A1 _07941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15334_ net1299 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12546_ net3240 net303 net404 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13159__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18053_ net1553 vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__buf_2
X_15265_ net1246 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12477_ net2533 net229 net412 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_4 _05490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12906__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17004_ clknet_leaf_134_wb_clk_i _02691_ _00987_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14216_ net1998 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11428_ _07679_ _07700_ team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1
+ vccd1 _07739_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_1663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15196_ net1174 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18038__1538 vssd1 vssd1 vccd1 vccd1 _18038__1538/HI net1538 sky130_fd_sc_hd__conb_1
XFILLER_0_26_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14147_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[39\] _04221_ _04233_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[71\]
+ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11359_ net1065 _07681_ vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__nand2_1
XANTENNA__10393__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09635__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14123__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14078_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[52\] _04236_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[124\]
+ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_60_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13029_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[57\] net2917 net866 vssd1 vssd1
+ vccd1 vccd1 _02096_ sky130_fd_sc_hd__mux2_1
X_17906_ net1426 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_59_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1060 team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1 vccd1
+ net1060 sky130_fd_sc_hd__buf_2
Xfanout1071 net1096 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__buf_2
XFILLER_0_20_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17837_ clknet_leaf_73_wb_clk_i net2420 _01777_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09550__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1082 net1089 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_2
Xfanout1093 net1095 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__buf_2
XFILLER_0_20_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08570_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[19\] net882 vssd1
+ vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__and3_1
X_17768_ clknet_leaf_85_wb_clk_i _03444_ _01708_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13634__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17967__1467 vssd1 vssd1 vccd1 vccd1 _17967__1467/HI net1467 sky130_fd_sc_hd__conb_1
XFILLER_0_18_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16719_ clknet_leaf_143_wb_clk_i _02406_ _00702_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17699_ clknet_leaf_101_wb_clk_i _03383_ _01640_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_117_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12000__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[14\] _04799_
+ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08714__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09053_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[12\] net908
+ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout212_A _07847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08433__B net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08004_ net1696 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[0\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09369__A2 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold510 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold521 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 team_01_WB.instance_to_wrap.cpu.c0.count\[13\] vssd1 vssd1 vccd1 vccd1 net2159
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12670__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold554 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[17\] vssd1 vssd1 vccd1 vccd1
+ net2170 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16201__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold565 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10384__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1121_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[58\] vssd1 vssd1 vccd1 vccd1
+ net2192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold587 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1219_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold598 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14114__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09955_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[3\] net974 vssd1
+ vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout679_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ net1105 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[2\] net927 vssd1
+ vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10136__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ net993 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[5\] net958 vssd1
+ vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__and3_1
Xhold1210 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[39\] vssd1 vssd1 vccd1 vccd1
+ net2837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1232 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2848 sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[1\] net671 net669 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__a22o_1
Xhold1243 team_01_WB.instance_to_wrap.cpu.K0.code\[4\] vssd1 vssd1 vccd1 vccd1 net2859
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout846_A net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1254 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1265 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[72\] vssd1 vssd1 vccd1 vccd1
+ net2881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2903 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09829__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[4\] net698 _05079_ _05083_
+ _05097_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__a2111o_1
Xhold1298 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[110\] vssd1 vssd1 vccd1 vccd1
+ net2914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10439__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08699_ _05030_ _05031_ _05037_ _05038_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__or4_2
XFILLER_0_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08501__B1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ _05115_ _07069_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10661_ _06438_ _06562_ net551 vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__mux2_1
XANTENNA__11034__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12845__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12400_ net2204 net203 net419 vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13380_ _03839_ _03840_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__nor2_1
X_10592_ net523 _06894_ _06906_ _06909_ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_1_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ net2595 net211 net430 vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15050_ net1272 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__inv_2
X_12262_ net2825 net218 net437 vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__mux2_1
XANTENNA__09158__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14001_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[9\] _04226_ _04254_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[97\]
+ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__a22o_1
X_11213_ net563 _07543_ _07544_ _07552_ vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__a31o_2
XFILLER_0_31_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12193_ net2883 net220 net445 vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__mux2_1
XANTENNA__12580__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10914__A2 _06526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14105__A2 _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ _07327_ _07329_ net535 vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__mux2_1
XANTENNA__09780__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_128_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__clkbuf_4
X_15952_ net1335 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__inv_2
X_11075_ _07413_ _07414_ _07359_ vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10026_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] _06365_ net623 vssd1
+ vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__mux2_2
X_14903_ net1195 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15883_ net1397 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__inv_2
XANTENNA__11924__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17622_ clknet_leaf_111_wb_clk_i _03307_ _01563_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_14834_ net1225 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13616__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17553_ clknet_leaf_17_wb_clk_i _03240_ _01536_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14765_ net1221 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__inv_2
X_11977_ net2965 net259 net473 vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__mux2_1
X_16504_ clknet_leaf_110_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[2\]
+ _00487_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13716_ _04103_ _04127_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[6\]
+ sky130_fd_sc_hd__nor2_1
X_10928_ net553 _07267_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__nor2_1
X_17484_ clknet_leaf_133_wb_clk_i _03171_ _01467_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14696_ net1346 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16435_ clknet_leaf_106_wb_clk_i _02189_ _00418_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13647_ net199 net196 _07925_ net645 vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__o211a_1
X_10859_ net375 _06707_ net372 _06671_ net533 net544 vssd1 vssd1 vccd1 vccd1 _07199_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_85_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13440__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16366_ clknet_leaf_69_wb_clk_i _02120_ _00349_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_13578_ _03914_ _03916_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18105_ net1590 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
X_15317_ net1219 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__inv_2
XANTENNA__16224__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12529_ net2269 net209 net405 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__mux2_1
X_16297_ clknet_leaf_59_wb_clk_i _02051_ _00280_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[20\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_26_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18036_ net1536 vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__buf_2
XFILLER_0_125_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15248_ net1272 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12355__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12490__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15179_ net1297 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10366__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16374__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 _07935_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_1
XANTENNA__09771__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout319 net321 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09740_ net1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[20\] net954
+ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__and3_1
XANTENNA__10118__B1 _04659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
.ends

