* NGSPICE file created from team_05.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt team_05 ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14] ADR_O[15]
+ ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22] ADR_O[23]
+ ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30] ADR_O[31]
+ ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0] DAT_I[10]
+ DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17] DAT_I[18]
+ DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25] DAT_I[26]
+ DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4] DAT_I[5]
+ DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12] DAT_O[13]
+ DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20] DAT_O[21]
+ DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28] DAT_O[29]
+ DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7] DAT_O[8]
+ DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O clk en gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5]
+ gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[0] gpio_oeb[10] gpio_oeb[11]
+ gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15] gpio_oeb[16] gpio_oeb[17] gpio_oeb[18]
+ gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21] gpio_oeb[22] gpio_oeb[23] gpio_oeb[24]
+ gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28] gpio_oeb[29] gpio_oeb[2] gpio_oeb[30]
+ gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7]
+ gpio_out[8] gpio_out[9] nrst vccd1 vssd1
XANTENNA__06501__B net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06883_ net311 _02438_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__nand2b_1
X_09671_ _03509_ _04102_ _04896_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08622_ _03913_ total_design.lcd_display.cnt_20ms\[4\] total_design.lcd_display.cnt_20ms\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__or3b_1
XANTENNA__11618__A0 _05630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ total_design.data_in_BUS\[12\] net342 _03900_ vssd1 vssd1 vccd1 vccd1 _03901_
+ sky130_fd_sc_hd__a21boi_1
XFILLER_0_77_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07504_ total_design.core.regFile.register\[14\]\[18\] net861 net853 total_design.core.regFile.register\[28\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08484_ _03813_ _03835_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__and2_1
XANTENNA__07837__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07435_ total_design.core.regFile.register\[29\]\[17\] net655 net562 total_design.core.regFile.register\[3\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09039__B2 _04290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout427_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12043__B1 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07366_ total_design.core.ctrl.instruction\[16\] _02846_ vssd1 vssd1 vccd1 vccd1
+ _02894_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_135_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11397__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06890__C total_design.core.ctrl.instruction\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_06317_ _01780_ _01804_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09105_ net325 _04170_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__nor2_1
XANTENNA__10185__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07297_ total_design.core.regFile.register\[14\]\[14\] net861 _01959_ total_design.core.regFile.register\[31\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__a22o_1
XANTENNA__08163__B _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_X net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09974__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09036_ _02113_ _04287_ net460 vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06248_ _01821_ _01825_ _01808_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout796_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold340 net49 vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
X_06179_ total_design.core.mem_ctrl.state\[1\] _01725_ vssd1 vssd1 vccd1 vccd1 _01761_
+ sky130_fd_sc_hd__nand2_1
Xhold351 net90 vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 total_design.lcd_display.row_2\[1\] vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold373 net55 vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 total_design.lcd_display.row_2\[48\] vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07222__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout963_A _01770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 total_design.lcd_display.row_2\[110\] vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout820 net822 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__buf_4
XANTENNA_fanout584_X net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout831 _01959_ vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_8
X_09938_ net207 net2161 net422 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__mux2_1
Xfanout842 net845 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_8
Xfanout853 _01949_ vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout864 _01943_ vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__buf_4
XANTENNA__06411__B net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout875 _01934_ vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__buf_8
XFILLER_0_99_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout886 _02023_ vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout897 net898 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_2
X_09869_ net211 net2432 net431 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__mux2_1
Xhold1040 total_design.core.regFile.register\[30\]\[31\] vssd1 vssd1 vccd1 vccd1 net2356
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 total_design.core.regFile.register\[24\]\[3\] vssd1 vssd1 vccd1 vccd1 net2367
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11900_ _05773_ _05774_ _05776_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__and3_1
Xhold1062 total_design.core.regFile.register\[22\]\[8\] vssd1 vssd1 vccd1 vccd1 net2378
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12880_ clknet_leaf_184_clk _00347_ net1037 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1073 total_design.core.regFile.register\[26\]\[5\] vssd1 vssd1 vccd1 vccd1 net2389
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 total_design.core.regFile.register\[10\]\[19\] vssd1 vssd1 vccd1 vccd1 net2400
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11609__A0 _05612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1095 total_design.core.regFile.register\[4\]\[7\] vssd1 vssd1 vccd1 vccd1 net2411
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07523__A total_design.core.ctrl.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ net1489 _05717_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_159_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14550_ net1270 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XANTENNA__07289__B1 _01986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11762_ net1817 net955 _05697_ _01880_ vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__a22o_1
XANTENNA__07828__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ clknet_leaf_14_clk _00968_ net1026 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10713_ net203 net2497 net359 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__mux2_1
X_14481_ clknet_leaf_33_clk _01548_ net1064 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_11693_ net28 net935 net878 net1842 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12034__B1 _05848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13432_ clknet_leaf_135_clk _00899_ net1187 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10644_ net218 net2286 net476 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13363_ clknet_leaf_178_clk _00830_ net1035 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10575_ net224 net2172 net372 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__mux2_1
XANTENNA__10095__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09884__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11986__Y _05848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12314_ total_design.core.math.pc_val\[19\] total_design.core.program_count.imm_val_reg\[19\]
+ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__and2_1
XANTENNA__07461__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13294_ clknet_leaf_190_clk _00761_ net1032 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12245_ net897 _02694_ _04541_ _05758_ _06088_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__o221a_1
XFILLER_0_121_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09185__A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ total_design.core.math.pc_val\[4\] total_design.core.program_count.imm_val_reg\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__nand2_1
XANTENNA__06567__A2 _01992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _05382_ _05383_ _05379_ _05381_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__a2bb2o_1
X_11058_ total_design.core.data_bus_o\[16\] net695 _05300_ net517 vssd1 vssd1 vccd1
+ vccd1 _05317_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11654__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ net195 net2504 net414 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__mux2_1
XANTENNA__10778__B total_design.core.data_bus_o\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09269__A1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11076__A1 total_design.core.data_bus_o\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14560__1280 vssd1 vssd1 vccd1 vccd1 _14560__1280/HI net1280 sky130_fd_sc_hd__conb_1
XANTENNA__10794__A _05049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07220_ total_design.core.regFile.register\[15\]\[13\] net607 net582 total_design.core.regFile.register\[6\]\[13\]
+ _02754_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_15_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12025__B1 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07151_ _02691_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10587__A0 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09794__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07082_ total_design.core.regFile.register\[24\]\[10\] net790 net786 total_design.core.regFile.register\[13\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__a22o_1
XANTENNA__07452__B1 _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14502__Q total_design.core.ctrl.instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout138 _05685_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout149 _05682_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__buf_4
X_07984_ total_design.core.regFile.register\[26\]\[28\] net870 net787 total_design.core.regFile.register\[13\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__a22o_1
X_09723_ net904 _04946_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__nor2_1
X_06935_ net551 net458 _02448_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11417__X _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11564__S net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09654_ net320 _04711_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_87_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06866_ total_design.core.regFile.register\[8\]\[6\] net804 _02419_ _02422_ vssd1
+ vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a211o_1
X_08605_ net1832 net339 net714 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[26\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_26_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06797_ total_design.core.regFile.register\[22\]\[5\] net676 net657 total_design.core.regFile.register\[29\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__a22o_1
X_09585_ _04730_ _04812_ net326 vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08158__B _02188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06730__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09969__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08468__C1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ total_design.keypad0.key_out\[13\] net932 _03843_ vssd1 vssd1 vccd1 vccd1
+ _03885_ sky130_fd_sc_hd__or3_1
XFILLER_0_132_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08467_ _03819_ _03820_ _03767_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12016__B1 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07418_ _02941_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__xnor2_4
X_08398_ _03752_ _03753_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__nor2_1
XANTENNA__07691__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08605__C net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07349_ total_design.core.regFile.register\[27\]\[15\] net781 _02878_ vssd1 vssd1
+ vccd1 vccd1 _02879_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_150_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06406__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06246__A1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10360_ net163 net2209 net489 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout799_X net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06797__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09276__Y _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ net472 _03369_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__nor2_1
X_10291_ net173 net2010 net498 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__mux2_1
XANTENNA__10643__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12030_ net123 net710 _05881_ _05890_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__o22a_1
XFILLER_0_131_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold170 total_design.core.instr_mem.instruction_adr_stored\[13\] vssd1 vssd1 vccd1
+ vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 total_design.lcd_display.lcd_rs vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold192 net50 vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_151_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout966_X net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout650 _02055_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout661 net662 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__buf_4
Xfanout672 net673 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__buf_4
X_13981_ clknet_leaf_92_clk _01161_ net1259 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[63\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout683 _02035_ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09499__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout694 _01933_ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11474__S net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12932_ clknet_leaf_105_clk _00399_ net1233 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_166_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14008__RESET_B net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12863_ clknet_leaf_183_clk _00330_ net1039 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06721__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11058__A1 total_design.core.data_bus_o\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09879__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11814_ net1881 _05707_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12794_ clknet_leaf_124_clk _00261_ net1186 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_164_Left_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09120__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ net1305 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_174_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ net1609 net958 net292 total_design.core.data_bus_o\[17\] vssd1 vssd1 vccd1
+ vccd1 _01373_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_174_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11073__A4 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12007__B1 _05810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14464_ clknet_leaf_52_clk net1446 net1094 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07682__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11676_ _05628_ net1610 net130 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__mux2_1
XANTENNA__13698__Q total_design.core.data_cpu_o\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07091__A_N _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13415_ clknet_leaf_19_clk _00882_ net1049 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10627_ net246 net1983 net476 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__mux2_1
X_14395_ net986 total_design.keypad0.next_rows\[1\] net1085 vssd1 vssd1 vccd1 vccd1
+ net113 sky130_fd_sc_hd__dfstp_1
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06316__B _01795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07434__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13346_ clknet_leaf_131_clk _00813_ net1197 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10558_ net161 net2647 net375 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11649__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10553__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13277_ clknet_leaf_10_clk _00744_ net1021 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10489_ net172 net1984 net378 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_173_Left_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12228_ net902 _02589_ _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12159_ total_design.core.math.pc_val\[2\] total_design.core.program_count.imm_val_reg\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10789__A total_design.core.data_bus_o\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06986__B _02515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06960__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ _02270_ _02282_ _02283_ _02284_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__or4_1
XANTENNA__12494__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06651_ total_design.core.regFile.register\[20\]\[2\] net671 net574 total_design.core.regFile.register\[24\]\[2\]
+ _02215_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a221o_1
XANTENNA__06712__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09789__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09370_ total_design.core.math.pc_val\[14\] _04583_ vssd1 vssd1 vccd1 vccd1 _04610_
+ sky130_fd_sc_hd__nor2_1
X_06582_ total_design.core.regFile.register\[22\]\[1\] net746 net735 net731 vssd1
+ vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_82_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire300_X net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08321_ total_design.core.data_mem.data_write_adr_reg\[18\] net546 net538 total_design.core.data_mem.data_read_adr_reg\[18\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07122__C1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11413__A _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08252_ net1372 net557 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[2\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_157_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07203_ _02718_ _02738_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__and2b_1
XFILLER_0_55_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08183_ net890 _03421_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[26\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07134_ total_design.core.regFile.register\[18\]\[11\] net857 net850 total_design.core.regFile.register\[9\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11772__A2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11559__S net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07065_ total_design.core.regFile.register\[27\]\[10\] net577 net566 total_design.core.regFile.register\[12\]\[10\]
+ _02609_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__a221o_1
XANTENNA__10463__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1034_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09029__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09717__A2 _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1201_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07967_ _03416_ _03420_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout661_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout759_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06951__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09706_ _03602_ net704 vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06918_ total_design.core.regFile.register\[18\]\[7\] net857 _01992_ total_design.core.regFile.register\[20\]\[7\]
+ _02471_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__a221o_1
XANTENNA__08169__A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ total_design.core.regFile.register\[30\]\[26\] net660 net602 total_design.core.regFile.register\[31\]\[26\]
+ _03397_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_104_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09637_ total_design.core.ctrl.instruction\[26\] net889 _04864_ net906 vssd1 vssd1
+ vccd1 vccd1 _04865_ sky130_fd_sc_hd__a22o_1
X_06849_ total_design.core.regFile.register\[29\]\[6\] net657 net568 total_design.core.regFile.register\[12\]\[6\]
+ _02405_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__a221o_1
XANTENNA__06703__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09568_ total_design.core.math.pc_val\[23\] _04777_ vssd1 vssd1 vccd1 vccd1 _04799_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_121_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08519_ _03868_ _03869_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10638__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ net297 _04357_ _04726_ _04732_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11460__A1 _05626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11530_ net1541 _05665_ net145 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11461_ net1550 _05677_ net155 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ clknet_leaf_184_clk _00667_ net1037 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10412_ net215 net1991 net385 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14180_ clknet_leaf_79_clk _01360_ net1218 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
X_11392_ net304 _05641_ _05610_ _05037_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_61_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11469__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13131_ clknet_leaf_114_clk _00598_ net1202 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10373__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10343_ net234 net2581 net491 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08351__B net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13062_ clknet_leaf_201_clk _00529_ net1004 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10274_ net242 net2550 net497 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12173__C1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ total_design.lcd_display.row_2\[57\] _05835_ _05847_ total_design.lcd_display.row_2\[33\]
+ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_167_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07195__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout480 _05011_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout491 _05006_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_4
X_13964_ clknet_leaf_111_clk _01144_ net1210 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09341__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ clknet_leaf_179_clk _00382_ net1034 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13895_ clknet_4_13__leaf_clk _01075_ net1221 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07352__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12846_ clknet_leaf_187_clk _00313_ net1028 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13895__RESET_B net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10548__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12777_ clknet_leaf_178_clk _00244_ net1032 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14516_ net1288 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XANTENNA__11451__A1 _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07655__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11728_ net73 net960 net293 net2690 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__a22o_1
XANTENNA__06327__A _01766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14447_ clknet_leaf_63_clk net1475 net1123 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ _05677_ net1706 net129 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07407__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14378_ clknet_leaf_4_clk _01519_ net1022 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold906 total_design.core.regFile.register\[4\]\[2\] vssd1 vssd1 vccd1 vccd1 net2222
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold917 total_design.core.regFile.register\[30\]\[5\] vssd1 vssd1 vccd1 vccd1 net2233
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13329_ clknet_leaf_148_clk _00796_ net1150 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10283__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold928 total_design.core.regFile.register\[12\]\[18\] vssd1 vssd1 vccd1 vccd1 net2244
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08080__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold939 total_design.core.regFile.register\[18\]\[23\] vssd1 vssd1 vccd1 vccd1 net2255
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08261__B net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_36_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08870_ net967 _04123_ _01921_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__o21a_4
XANTENNA__07186__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07821_ _03323_ _03325_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06933__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ total_design.core.regFile.register\[23\]\[23\] net678 net674 total_design.core.regFile.register\[22\]\[23\]
+ _03255_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_84_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06703_ total_design.core.regFile.register\[20\]\[3\] net670 net581 total_design.core.regFile.register\[6\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a22o_1
X_07683_ total_design.core.regFile.register\[16\]\[22\] net855 net847 total_design.core.regFile.register\[15\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__a22o_1
X_09422_ _04638_ _04658_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__nor2_1
XANTENNA__12219__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06634_ total_design.core.regFile.register\[20\]\[2\] net818 net815 total_design.core.regFile.register\[4\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__a22o_1
XANTENNA__07621__A _03112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ _02841_ _04568_ _04591_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__or3_1
XFILLER_0_158_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10458__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06565_ total_design.core.regFile.register\[21\]\[1\] net759 _02119_ _02121_ _02127_
+ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08304_ net1466 net940 _03686_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[9\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11442__A1 _05636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06496_ net741 net733 net724 vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__and3_1
X_09284_ _04482_ _04526_ net463 vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07110__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11993__A2 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08235_ net1482 net542 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[18\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_160_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1151_A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout507_A _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09548__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08166_ net892 _02589_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[9\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07117_ total_design.core.regFile.register\[13\]\[11\] net669 net639 total_design.core.regFile.register\[2\]\[11\]
+ _02658_ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__a221o_1
X_08097_ total_design.core.regFile.register\[7\]\[30\] net654 net635 total_design.core.regFile.register\[16\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__a22o_1
XANTENNA__08071__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10193__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08171__B _02845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09982__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload90 clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 clkload90/Y sky130_fd_sc_hd__clkinv_4
X_07048_ _02593_ vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[10\] sky130_fd_sc_hd__inv_2
XANTENNA_fanout876_A _01934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07177__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _04249_ _04251_ net468 vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__mux2_1
XANTENNA__06924__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_162_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10961_ total_design.core.data_bus_o\[3\] net697 vssd1 vssd1 vccd1 vccd1 _05220_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_X net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ clknet_leaf_30_clk _00167_ net1060 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13680_ clknet_leaf_48_clk total_design.core.data_mem.data_read_adr_i\[20\] net1102
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[20\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07885__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10892_ _05135_ _05139_ _05137_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a21oi_2
X_12631_ clknet_leaf_123_clk _00098_ net1166 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10368__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12562_ net1419 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07101__A2 total_design.core.ctrl.instruction\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14301_ clknet_leaf_103_clk _00015_ net1239 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11513_ net1529 _05643_ net150 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12493_ net977 total_design.core.instr_mem.instruction_i\[10\] vssd1 vssd1 vccd1
+ vccd1 _01701_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14232_ clknet_leaf_60_clk _01412_ net1132 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dfrtp_1
X_11444_ net1565 _05612_ net157 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14163_ clknet_leaf_34_clk _01343_ net1066 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11375_ _05627_ _05631_ _05632_ _05633_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__and4_1
XFILLER_0_1_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09892__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13114_ clknet_leaf_132_clk _00581_ net1196 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10326_ net165 net2578 net494 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__mux2_1
X_14094_ clknet_leaf_101_clk _01274_ net1237 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06313__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_2__f_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_13045_ clknet_leaf_167_clk _00512_ net1155 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10257_ net176 net2024 net501 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1220 net1221 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07168__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1231 net1232 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__clkbuf_2
Xfanout1242 net1243 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__clkbuf_2
X_10188_ net286 net2475 net390 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__mux2_1
Xfanout1253 net1257 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__clkbuf_4
Xfanout1264 net1265 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__buf_2
XANTENNA__06915__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13947_ clknet_leaf_89_clk _01127_ net1260 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11662__S net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07876__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ clknet_leaf_26_clk total_design.core.ctrl.imm_32\[17\] net1107 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07340__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12829_ clknet_leaf_9_clk _00296_ net1020 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10278__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09078__C1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08256__B net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06350_ _01917_ _01920_ _01739_ _01915_ vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__a211o_1
XANTENNA__11424__A1 _05358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07628__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06281_ total_design.core.instr_mem.instruction_adr_i\[4\] total_design.core.instr_mem.instruction_adr_stored\[4\]
+ net984 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_150_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_150_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08020_ total_design.core.regFile.register\[14\]\[29\] net861 net759 total_design.core.regFile.register\[21\]\[29\]
+ _03515_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold703 total_design.core.regFile.register\[7\]\[6\] vssd1 vssd1 vccd1 vccd1 net2019
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11410__B _05064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold714 total_design.core.regFile.register\[5\]\[13\] vssd1 vssd1 vccd1 vccd1 net2030
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold725 total_design.core.regFile.register\[31\]\[11\] vssd1 vssd1 vccd1 vccd1 net2041
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 total_design.core.regFile.register\[3\]\[31\] vssd1 vssd1 vccd1 vccd1 net2052
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 total_design.core.regFile.register\[17\]\[9\] vssd1 vssd1 vccd1 vccd1 net2063
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold758 total_design.core.regFile.register\[4\]\[15\] vssd1 vssd1 vccd1 vccd1 net2074
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07800__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09971_ net211 net2414 net419 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__mux2_1
Xhold769 total_design.core.regFile.register\[27\]\[12\] vssd1 vssd1 vccd1 vccd1 net2085
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08922_ net473 _03112_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12152__A2 _05832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08853_ _04107_ _04104_ _04074_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1403 total_design.core.regFile.register\[1\]\[17\] vssd1 vssd1 vccd1 vccd1 net2719
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout192_A _04822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1414 total_design.core.regFile.register\[19\]\[14\] vssd1 vssd1 vccd1 vccd1 net2730
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1425 total_design.core.regFile.register\[4\]\[17\] vssd1 vssd1 vccd1 vccd1 net2741
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06906__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1436 total_design.core.regFile.register\[28\]\[31\] vssd1 vssd1 vccd1 vccd1 net2752
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07804_ total_design.core.regFile.register\[11\]\[24\] net613 net574 total_design.core.regFile.register\[24\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1447 total_design.core.regFile.register\[6\]\[6\] vssd1 vssd1 vccd1 vccd1 net2763
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08784_ _02613_ net310 vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__and2_1
Xhold1458 total_design.core.regFile.register\[21\]\[6\] vssd1 vssd1 vccd1 vccd1 net2774
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1469 total_design.core.data_bus_o\[19\] vssd1 vssd1 vccd1 vccd1 net2785 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_140_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07735_ total_design.core.regFile.register\[26\]\[23\] net869 net798 total_design.core.regFile.register\[29\]\[23\]
+ _03238_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_140_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11572__S net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1199_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07867__B1 total_design.core.ctrl.imm_32\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09550__B _04776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07666_ total_design.core.regFile.register\[0\]\[21\] net684 _03159_ _03176_ vssd1
+ vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_149_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07331__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09405_ _02941_ _04102_ _04184_ _04191_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__a22oi_1
X_06617_ _02116_ _02187_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__xnor2_4
XANTENNA__09069__C1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10188__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07597_ _03096_ _03099_ _03100_ _03110_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout624_A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09977__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07619__B1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09336_ net318 _04382_ _04576_ net295 vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__a211o_1
X_06548_ total_design.core.regFile.register\[31\]\[1\] net925 net911 net946 vssd1
+ vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__and4_1
XFILLER_0_164_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11966__A2 _05826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ _02637_ net508 net504 _02635_ _04510_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_141_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_141_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06479_ total_design.core.regFile.register\[29\]\[0\] net747 net729 net727 vssd1
+ vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout1154_X net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08218_ net1429 net544 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[1\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09278__A _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09198_ _02489_ net447 net289 _04443_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout993_A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08149_ total_design.core.regFile.register\[22\]\[31\] net675 net605 total_design.core.regFile.register\[15\]\[31\]
+ _03625_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__a221o_1
XANTENNA__08044__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06414__B net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07398__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11160_ _05418_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10111_ net191 net2802 net404 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11091_ _05057_ _05266_ _05267_ _05278_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__a31o_1
XANTENNA__10651__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12143__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09544__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10042_ net199 net2618 net411 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__mux2_1
Xhold30 total_design.core.data_mem.data_read_adr_reg\[21\] vssd1 vssd1 vccd1 vccd1
+ net1346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 total_design.core.data_mem.data_cpu_i_reg\[30\] vssd1 vssd1 vccd1 vccd1 net1357
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 total_design.core.data_mem.data_bus_i_reg\[4\] vssd1 vssd1 vccd1 vccd1 net1368
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 total_design.core.math.pc_val\[23\] vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold74 total_design.core.data_mem.data_cpu_i_reg\[8\] vssd1 vssd1 vccd1 vccd1 net1390
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 total_design.core.data_mem.data_cpu_i_reg\[25\] vssd1 vssd1 vccd1 vccd1 net1401
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 total_design.core.instr_mem.instruction_adr_stored\[31\] vssd1 vssd1 vccd1
+ vccd1 net1412 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ clknet_leaf_76_clk total_design.core.data_mem.data_cpu_i\[10\] net1213 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[10\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11103__B1 _05361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ total_design.lcd_display.row_2\[80\] _05818_ _05840_ total_design.lcd_display.row_1\[48\]
+ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__a22o_1
XANTENNA__11482__S net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13732_ clknet_leaf_76_clk total_design.core.data_mem.stored_write_data\[7\] net1213
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[7\] sky130_fd_sc_hd__dfrtp_2
Xclkbuf_4_10__f_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10944_ _05178_ _05200_ _05202_ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__a21boi_2
XANTENNA__07858__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07322__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13663_ clknet_leaf_61_clk total_design.core.data_mem.data_read_adr_i\[3\] net1129
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10098__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10875_ _01885_ _05133_ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09887__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12614_ clknet_leaf_198_clk _00081_ net1001 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13594_ clknet_leaf_34_clk total_design.core.data_mem.data_bus_i\[30\] net1067 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12545_ net1387 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_132_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_132_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_164_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12476_ net980 net2476 net884 _01692_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14215_ clknet_leaf_78_clk _01395_ net1217 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfrtp_1
X_11427_ net1552 _05663_ net157 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__mux2_1
XANTENNA_5 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06324__B _01900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09783__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14146_ clknet_leaf_43_clk _01326_ net1083 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output86_A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14204__RESET_B net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11358_ _05459_ _05475_ _05616_ _05471_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11590__A0 _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11657__S net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ net230 net1955 net495 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__mux2_1
XANTENNA__10561__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14077_ clknet_leaf_85_clk _01257_ net1258 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[95\]
+ sky130_fd_sc_hd__dfrtp_1
X_11289_ _05543_ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_5_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13028_ clknet_leaf_108_clk _00495_ net1224 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_199_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_199_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06349__B1 total_design.core.ctrl.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_174_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1050 net1051 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_4
Xfanout1061 net1065 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__clkbuf_4
Xfanout1072 net1081 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__clkbuf_4
Xfanout1083 net1084 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08819__X _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1094 net1095 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07561__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09651__A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07520_ _03038_ _03039_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07849__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06339__X _01915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07451_ total_design.core.regFile.register\[23\]\[17\] net810 net759 total_design.core.regFile.register\[21\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09797__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06402_ net923 net914 net912 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__and3_1
X_07382_ total_design.core.regFile.register\[2\]\[16\] net638 net622 total_design.core.regFile.register\[4\]\[16\]
+ _02908_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__a221o_1
XANTENNA__09066__A2 _04283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09121_ total_design.core.math.pc_val\[2\] total_design.core.math.pc_val\[3\] total_design.core.math.pc_val\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_44_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06333_ wishbone.curr_state\[2\] wishbone.curr_state\[1\] vssd1 vssd1 vccd1 vccd1
+ _01912_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_123_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06264_ _01771_ _01842_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__nor2_1
X_09052_ _04181_ _04131_ net459 vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08003_ total_design.core.regFile.register\[9\]\[28\] net665 net622 total_design.core.regFile.register\[4\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__a22o_1
XANTENNA__08026__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06195_ total_design.core.mem_ctrl.state\[1\] total_design.core.mem_ctrl.state\[0\]
+ total_design.core.mem_ctrl.state\[2\] vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__or3b_1
XFILLER_0_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold500 total_design.lcd_display.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 net46 vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 net47 vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout205_A _04740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold533 total_design.lcd_display.row_1\[61\] vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09774__A0 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold544 total_design.core.regFile.register\[12\]\[0\] vssd1 vssd1 vccd1 vccd1 net1860
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08730__A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11581__A0 _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold555 total_design.lcd_display.cnt_20ms\[3\] vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 total_design.data_in_BUS\[10\] vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11567__S net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold577 total_design.core.regFile.register\[27\]\[0\] vssd1 vssd1 vccd1 vccd1 net1893
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 total_design.core.regFile.register\[31\]\[27\] vssd1 vssd1 vccd1 vccd1 net1904
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07617__Y _03131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10471__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09954_ net278 net2166 net419 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__mux2_1
Xhold599 total_design.core.regFile.register\[2\]\[2\] vssd1 vssd1 vccd1 vccd1 net1915
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12125__A2 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08905_ _02338_ _04098_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__nand2_2
XFILLER_0_148_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06250__A _01771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09885_ net244 net2482 net426 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout574_A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1200 total_design.core.regFile.register\[26\]\[11\] vssd1 vssd1 vccd1 vccd1 net2516
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 total_design.core.regFile.register\[4\]\[16\] vssd1 vssd1 vccd1 vccd1 net2527
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1222 total_design.core.regFile.register\[25\]\[23\] vssd1 vssd1 vccd1 vccd1 net2538
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ _04006_ _04009_ _04010_ _04002_ _04000_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__o221a_1
Xhold1233 total_design.core.regFile.register\[27\]\[2\] vssd1 vssd1 vccd1 vccd1 net2549
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 total_design.core.regFile.register\[5\]\[3\] vssd1 vssd1 vccd1 vccd1 net2560
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1255 total_design.core.regFile.register\[2\]\[14\] vssd1 vssd1 vccd1 vccd1 net2571
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 total_design.core.regFile.register\[27\]\[22\] vssd1 vssd1 vccd1 vccd1 net2582
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07552__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1277 total_design.core.regFile.register\[18\]\[31\] vssd1 vssd1 vccd1 vccd1 net2593
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ _04021_ _04017_ _04019_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__and3b_1
XANTENNA__06760__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1288 total_design.core.regFile.register\[10\]\[8\] vssd1 vssd1 vccd1 vccd1 net2604
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1299 total_design.core.regFile.register\[19\]\[16\] vssd1 vssd1 vccd1 vccd1 net2615
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout839_A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07718_ _03207_ _03226_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_68_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ net1819 _03954_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_68_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07649_ total_design.core.regFile.register\[22\]\[21\] net675 net667 total_design.core.regFile.register\[13\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06409__B net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10660_ net244 net1885 net364 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06542__A_N _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09319_ total_design.core.math.pc_val\[12\] _04539_ vssd1 vssd1 vccd1 vccd1 _04561_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10646__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10591_ net161 net2791 net371 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_114_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12330_ total_design.core.math.pc_val\[21\] total_design.core.program_count.imm_val_reg\[21\]
+ vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__and2_1
XANTENNA__12809__RESET_B net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout996_X net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08017__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ net996 _04585_ net895 vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14000_ clknet_leaf_83_clk _01180_ net1241 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11212_ _05456_ net294 _05467_ _05469_ _05356_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__o32ai_4
X_12192_ net898 _06041_ net526 vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11572__A0 _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11477__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__clkbuf_4
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__clkbuf_4
X_11143_ _05390_ _05394_ _05400_ _05393_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__o22ai_1
XANTENNA__10381__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12116__A2 _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07791__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XANTENNA__07256__A _02770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
X_11074_ net518 _05059_ _05134_ _05044_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__o211a_1
XANTENNA__06160__A total_design.core.ctrl.instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10025_ net259 net2083 net412 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__mux2_1
XANTENNA__07543__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output124_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11088__C1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11976_ _05811_ _05820_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__nor2_4
X_13715_ clknet_leaf_27_clk total_design.core.data_mem.stored_read_data\[22\] net1077
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[22\] sky130_fd_sc_hd__dfrtp_1
X_10927_ _05155_ _05157_ _05159_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13646_ clknet_leaf_49_clk total_design.core.data_mem.data_write_adr_i\[18\] net1101
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[18\] sky130_fd_sc_hd__dfrtp_1
X_10858_ _05116_ _05096_ _05092_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13577_ clknet_leaf_35_clk total_design.core.data_mem.data_bus_i\[13\] net1071 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[13\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10556__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_105_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10789_ total_design.core.data_bus_o\[7\] net698 vssd1 vssd1 vccd1 vccd1 _05048_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12528_ net978 total_design.core.ctrl.instruction\[27\] net883 _01718_ vssd1 vssd1
+ vccd1 vccd1 _01566_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12459_ net2103 net172 net346 vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14129_ clknet_leaf_96_clk _01309_ net1253 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10291__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12107__A2 _05812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07782__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ total_design.core.regFile.register\[25\]\[8\] net649 net630 total_design.core.regFile.register\[5\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06501__C net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _03508_ net505 _04188_ _03507_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__a2bb2o_1
X_06882_ net555 total_design.core.data_mem.data_cpu_i\[6\] total_design.core.ctrl.imm_32\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07534__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08621_ total_design.lcd_display.cnt_20ms\[9\] total_design.lcd_display.cnt_20ms\[8\]
+ total_design.lcd_display.cnt_20ms\[7\] total_design.lcd_display.cnt_20ms\[6\] vssd1
+ vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__or4bb_1
XANTENNA__06742__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08552_ _03889_ _03893_ _03898_ _03899_ _03767_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__a311o_1
XFILLER_0_89_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07503_ total_design.core.regFile.register\[12\]\[18\] _01980_ net758 total_design.core.regFile.register\[4\]\[18\]
+ _03023_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_46_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08483_ _03813_ _03835_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__nor2_1
XANTENNA__12291__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout155_A _05681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07434_ total_design.core.regFile.register\[7\]\[17\] net651 net608 total_design.core.regFile.register\[18\]\[17\]
+ _02957_ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__a221o_1
XANTENNA__09039__A2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07365_ net751 _02893_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[15\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10466__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12247__A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout322_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09104_ net326 _04165_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__nand2_1
X_06316_ _01784_ _01795_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_33_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07296_ total_design.core.regFile.register\[7\]\[14\] net770 _02828_ vssd1 vssd1
+ vccd1 vccd1 _02829_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09035_ _04150_ _04153_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__or2_1
X_06247_ _01808_ _01825_ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold330 total_design.lcd_display.row_2\[51\] vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06178_ total_design.core.mem_ctrl.state\[0\] total_design.core.mem_ctrl.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__nand2_1
Xhold341 total_design.lcd_display.row_1\[83\] vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11554__A0 _05477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold352 total_design.lcd_display.row_2\[55\] vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09211__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout691_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 total_design.data_in_BUS\[9\] vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 total_design.lcd_display.row_2\[42\] vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold385 total_design.lcd_display.row_2\[65\] vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 total_design.lcd_display.row_2\[56\] vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09990__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout810 net813 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_8
Xfanout821 net822 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__buf_4
X_09937_ net211 net2557 net423 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__mux2_1
Xfanout832 net833 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__buf_4
Xfanout843 net845 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10214__B net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout956_A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_X net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 _01947_ vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06411__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout865 _01941_ vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout876 _01934_ vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__buf_4
Xfanout887 _02023_ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_2
X_09868_ net216 net2091 net430 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__mux2_1
Xfanout898 _02017_ vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__buf_2
Xhold1030 total_design.core.regFile.register\[9\]\[17\] vssd1 vssd1 vccd1 vccd1 net2346
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 total_design.core.regFile.register\[28\]\[25\] vssd1 vssd1 vccd1 vccd1 net2357
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 total_design.core.regFile.register\[4\]\[23\] vssd1 vssd1 vccd1 vccd1 net2368
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ _04033_ _04057_ _04063_ _04073_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__or4_2
Xhold1063 total_design.core.regFile.register\[6\]\[4\] vssd1 vssd1 vccd1 vccd1 net2379
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 total_design.core.regFile.register\[9\]\[25\] vssd1 vssd1 vccd1 vccd1 net2390
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06733__B1 _01992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09799_ net216 net2614 net438 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__mux2_1
Xhold1085 total_design.core.regFile.register\[19\]\[20\] vssd1 vssd1 vccd1 vccd1 net2401
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1096 total_design.core.regFile.register\[29\]\[15\] vssd1 vssd1 vccd1 vccd1 net2412
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ _05717_ _05718_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_107_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ net1823 net955 _05697_ _01876_ vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09683__C1 _04904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13500_ clknet_leaf_30_clk _00967_ net1060 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10712_ net205 net2308 net357 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14480_ clknet_leaf_38_clk _01547_ net1079 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_11692_ net27 net937 _05690_ net2671 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_3__f_clk_X clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09230__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13431_ clknet_leaf_124_clk _00898_ net1186 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10643_ net214 net2287 net476 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10376__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10229__X _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09986__A0 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13362_ clknet_leaf_139_clk _00829_ net1185 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_172_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10574_ net234 net2474 net369 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__mux2_1
XANTENNA__06155__A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11793__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12313_ total_design.core.math.pc_val\[19\] total_design.core.program_count.imm_val_reg\[19\]
+ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13293_ clknet_leaf_0_clk _00760_ net1005 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12337__A2 _03187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12244_ _06086_ _06087_ _05760_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__or3b_1
XFILLER_0_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06438__A_N total_design.core.ctrl.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12175_ _06026_ total_design.core.math.pc_val\[3\] net526 vssd1 vssd1 vccd1 vccd1
+ _01473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07764__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ _05384_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__inv_2
XANTENNA__06972__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ _05243_ _05304_ _05295_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_64_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10008_ net200 net2770 net416 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_95_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10778__C _05028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11076__A2 total_design.core.data_bus_o\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11959_ _05798_ _05820_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__nor2_4
XFILLER_0_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14547__A total_design.lcd_display.lcd_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11670__S net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13629_ clknet_leaf_62_clk total_design.core.data_mem.data_write_adr_i\[1\] net1128
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10286__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09426__C1 _04105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08264__B net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07150_ _02666_ _02687_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07081_ total_design.core.regFile.register\[20\]\[10\] _01992_ net758 total_design.core.regFile.register\[4\]\[10\]
+ _02615_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_130_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06660__C1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06512__B net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07755__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout139 _05685_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_4
X_07983_ total_design.core.regFile.register\[25\]\[28\] net843 net765 total_design.core.regFile.register\[6\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_4_14__f_clk_X clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ _04944_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__nand2b_1
X_06934_ net458 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[7\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_129_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09901__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12500__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09653_ net329 _04793_ _04878_ net319 vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06865_ total_design.core.regFile.register\[10\]\[6\] net835 _02420_ _02421_ vssd1
+ vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08604_ net2884 net338 net714 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[25\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_171_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09584_ _03326_ net509 net296 _04466_ _04813_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_26_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06796_ total_design.core.regFile.register\[23\]\[5\] net680 _02355_ net688 vssd1
+ vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_26_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08535_ net717 _03884_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[10\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout158_X net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11580__S net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1181_A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout537_A _04100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11433__X _05679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08466_ _03791_ _03794_ _03818_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__nand3_1
XFILLER_0_37_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07140__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__Y _05411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07417_ _02890_ _02942_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_154_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08397_ _03751_ total_design.keypad0.key_out\[4\] total_design.keypad0.key_out\[6\]
+ _03714_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout704_A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08174__B _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07348_ total_design.core.regFile.register\[9\]\[15\] net852 net829 total_design.core.regFile.register\[1\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11775__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07279_ total_design.core.regFile.register\[11\]\[14\] net615 net588 total_design.core.regFile.register\[28\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12319__A2 _03090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07994__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09018_ net335 _03415_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10290_ net178 net1912 net498 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold160 total_design.key_data vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 total_design.core.data_mem.data_read_adr_reg2\[28\] vssd1 vssd1 vccd1 vccd1
+ net1487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 total_design.core.data_mem.data_read_adr_reg2\[13\] vssd1 vssd1 vccd1 vccd1
+ net1498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 total_design.data_in_BUS\[11\] vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09573__X _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_X net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 net643 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_109_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout651 _02054_ vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_109_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout662 _02050_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__buf_4
X_13980_ clknet_leaf_109_clk _01160_ net1228 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[62\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout673 _02042_ vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__buf_4
Xfanout684 _02035_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_6
Xfanout695 net696 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__buf_2
X_12931_ clknet_leaf_15_clk _00398_ net1022 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06706__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07903__C1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12862_ clknet_leaf_157_clk _00329_ net1141 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11813_ total_design.lcd_display.cnt_20ms\[9\] _05707_ vssd1 vssd1 vccd1 vccd1 _05709_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10895__A total_design.core.data_bus_o\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12793_ clknet_leaf_195_clk _00260_ net1010 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11490__S net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14532_ net1304 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XFILLER_0_84_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ net1621 net959 net292 total_design.core.data_bus_o\[16\] vssd1 vssd1 vccd1
+ vccd1 _01372_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07131__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09671__A2 _04102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14463_ clknet_leaf_51_clk net1867 net1093 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11675_ _05612_ net1709 net129 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13414_ clknet_leaf_200_clk _00881_ net1004 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09895__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10626_ net287 net2494 net479 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__mux2_1
X_14394_ net986 total_design.keypad0.next_rows\[0\] net1085 vssd1 vssd1 vccd1 vccd1
+ net112 sky130_fd_sc_hd__dfrtp_1
X_13345_ clknet_leaf_118_clk _00812_ net1169 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10557_ net167 total_design.core.regFile.register\[6\]\[30\] net376 vssd1 vssd1 vccd1
+ vccd1 _00837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07985__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13276_ clknet_leaf_10_clk _00743_ net1020 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10488_ net179 net2179 net378 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__mux2_1
X_12227_ _04494_ _05757_ _05760_ _06072_ net527 vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ net1497 _03928_ _06011_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__a21o_1
XANTENNA__11665__S net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ _05360_ _05363_ _05364_ _05366_ _05367_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__o32ai_4
XANTENNA__08781__A_N total_design.core.data_mem.data_cpu_i\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12089_ total_design.lcd_display.row_1\[100\] _05810_ _05850_ total_design.lcd_display.row_2\[4\]
+ _05946_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_34_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08259__B net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06650_ total_design.core.regFile.register\[16\]\[2\] net632 net628 total_design.core.regFile.register\[5\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06581_ total_design.core.regFile.register\[0\]\[1\] net683 vssd1 vssd1 vccd1 vccd1
+ _02152_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_82_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09111__A1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08320_ net1494 net939 _03694_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[17\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11413__B _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08251_ net1417 net557 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[1\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06507__B net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07202_ _02739_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08182_ net890 _03375_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[25\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11757__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07133_ total_design.core.regFile.register\[30\]\[11\] net841 net809 total_design.core.regFile.register\[5\]\[11\]
+ _02674_ vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07976__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07064_ total_design.core.regFile.register\[25\]\[10\] net647 net589 total_design.core.regFile.register\[1\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07728__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1027_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__A1 _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11575__S net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout487_A _05007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07625__Y _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09553__B _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ _03462_ _03464_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__and2_2
X_09705_ net169 net2489 net453 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06917_ total_design.core.regFile.register\[24\]\[7\] net790 net783 total_design.core.regFile.register\[2\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__a22o_1
X_07897_ total_design.core.regFile.register\[19\]\[26\] net641 net609 total_design.core.regFile.register\[18\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__a22o_1
XANTENNA__08169__B _02746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout654_A _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09636_ _04863_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06848_ total_design.core.regFile.register\[26\]\[6\] net645 net591 total_design.core.regFile.register\[1\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07900__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09567_ net449 _04797_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06779_ _02339_ _02340_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08518_ _03852_ _03867_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__and2_1
XANTENNA__07113__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09498_ _04551_ _04687_ _04731_ net289 _04728_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__o221a_1
XFILLER_0_136_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11996__B1 _05829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08449_ net931 _01759_ _03800_ _03801_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__or4_1
XFILLER_0_81_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11460_ net1535 _05626_ net156 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_5_0_clk_X clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09405__A2 _04102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10411_ net223 net1890 net387 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__mux2_1
X_11391_ total_design.core.data_bus_o\[29\] net697 net303 _05641_ net510 vssd1 vssd1
+ vccd1 vccd1 _05650_ sky130_fd_sc_hd__a221o_4
XANTENNA__10654__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13130_ clknet_leaf_22_clk _00597_ net1049 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10342_ net229 net2714 net488 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08351__C _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13061_ clknet_leaf_116_clk _00528_ net1203 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10273_ net256 net2341 net496 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12012_ total_design.lcd_display.row_1\[81\] _05815_ _05827_ total_design.lcd_display.row_1\[33\]
+ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__a22o_1
XANTENNA__09744__A _04121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06927__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11485__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08392__A2 _01905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout470 _02111_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_4
Xfanout481 _05011_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout492 net495 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__buf_6
X_13963_ clknet_leaf_93_clk _01143_ net1255 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_85_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12914_ clknet_leaf_145_clk _00381_ net1177 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13894_ clknet_leaf_73_clk _01074_ net1209 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07352__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12228__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ clknet_leaf_2_clk _00312_ net1014 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12776_ clknet_leaf_23_clk _00243_ net1055 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08301__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11727_ net699 _05695_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__and2_1
X_14515_ net1287 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_72_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08852__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11658_ _05626_ net1774 net131 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__mux2_1
X_14446_ clknet_leaf_63_clk net1355 net1130 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10609_ net222 net2527 net367 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__mux2_1
XANTENNA__10564__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14377_ clknet_leaf_174_clk _01518_ net1156 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11589_ _05618_ net1741 net137 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10791__C total_design.core.data_bus_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07958__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold907 total_design.core.data_bus_o\[2\] vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold918 total_design.core.regFile.register\[17\]\[19\] vssd1 vssd1 vccd1 vccd1 net2234
+ sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ clknet_leaf_184_clk _00795_ net1039 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold929 total_design.core.regFile.register\[28\]\[13\] vssd1 vssd1 vccd1 vccd1 net2245
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06630__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13259_ clknet_leaf_120_clk _00726_ net1171 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06918__B1 _01992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07820_ _03324_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07591__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ total_design.core.regFile.register\[5\]\[23\] net628 net581 total_design.core.regFile.register\[6\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_76_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06702_ _02213_ _02239_ _02238_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08135__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07682_ total_design.core.regFile.register\[9\]\[22\] net851 net795 total_design.core.regFile.register\[11\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__a22o_1
XANTENNA__07343__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09421_ _02918_ _02937_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__nor2_1
XANTENNA__12219__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06633_ _02189_ _02200_ _02201_ _02202_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__or4_1
XFILLER_0_149_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09352_ _04568_ _04591_ _02841_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09096__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06564_ total_design.core.regFile.register\[7\]\[1\] net920 net911 net907 vssd1 vssd1
+ vccd1 vccd1 _02137_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08303_ total_design.core.data_mem.data_write_adr_reg\[9\] net548 net540 total_design.core.data_mem.data_read_adr_reg\[9\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_150_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09283_ _04225_ _04228_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__nand2_1
X_06495_ total_design.core.regFile.register\[10\]\[0\] net740 net731 net723 vssd1
+ vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08234_ net1450 net542 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[17\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_51_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__A _02188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08165_ _02021_ _02540_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[8\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__10474__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout402_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1144_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07116_ total_design.core.regFile.register\[18\]\[11\] net611 net565 total_design.core.regFile.register\[3\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__a22o_1
XANTENNA__07949__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_165_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08096_ total_design.core.regFile.register\[22\]\[30\] net676 net614 total_design.core.regFile.register\[11\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload80 clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__inv_6
Xclkload91 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 clkload91/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06621__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07047_ net721 _02590_ _02591_ _02592_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout771_A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06909__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08998_ net335 net299 _04250_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__a21o_1
XANTENNA__07582__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ total_design.core.regFile.register\[26\]\[27\] net645 net575 total_design.core.regFile.register\[24\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_3_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_67_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08126__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_170_Right_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ _05188_ _05190_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ _04845_ _04846_ net704 vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06688__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ _05149_ _05147_ _05104_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__mux2_1
XANTENNA__10649__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12630_ clknet_leaf_153_clk _00097_ net1138 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12561_ net1437 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11512_ net1579 _05648_ net152 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14300_ clknet_leaf_103_clk _00014_ net1239 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12492_ net975 total_design.core.ctrl.instruction\[9\] net881 _01700_ vssd1 vssd1
+ vccd1 vccd1 _01548_ sky130_fd_sc_hd__a22o_1
X_14231_ clknet_leaf_56_clk _01411_ net1115 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dfrtp_1
X_11443_ net1613 _05609_ net160 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__mux2_1
XANTENNA__10384__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14162_ clknet_leaf_31_clk _01342_ net1060 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11374_ total_design.core.data_bus_o\[28\] net700 _05610_ vssd1 vssd1 vccd1 vccd1
+ _05633_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_169_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13113_ clknet_leaf_188_clk _00580_ net1028 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10325_ net169 net2267 net492 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__mux2_1
X_14093_ clknet_leaf_89_clk _01273_ net1258 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12146__B1 _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13044_ clknet_leaf_144_clk _00511_ net1176 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07546__X _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10256_ net182 net2442 net501 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__mux2_1
XANTENNA__06450__X total_design.core.ctrl.imm_32\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1210 net1211 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__clkbuf_2
Xfanout1221 net1222 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__buf_4
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1232 net1240 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__clkbuf_2
X_10187_ _04116_ _04120_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__or2_1
Xfanout1243 net1252 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1254 net1257 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__clkbuf_4
Xfanout1265 net39 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_58_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08117__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13946_ clknet_leaf_86_clk _01126_ net1248 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07325__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06679__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13877_ clknet_leaf_26_clk total_design.core.ctrl.imm_32\[16\] net1107 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[16\] sky130_fd_sc_hd__dfrtp_1
X_12828_ clknet_leaf_30_clk _00295_ net1064 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12759_ clknet_leaf_162_clk _00226_ net1166 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_max_cap288_X net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06280_ net930 _01854_ _01857_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10294__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06851__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14429_ clknet_leaf_33_clk total_design.core.data_out_INSTR\[24\] net1070 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold704 total_design.core.regFile.register\[19\]\[29\] vssd1 vssd1 vccd1 vccd1 net2020
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 total_design.data_in_BUS\[5\] vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
Xwire690 _02009_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold726 total_design.core.regFile.register\[23\]\[3\] vssd1 vssd1 vccd1 vccd1 net2042
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold737 total_design.core.regFile.register\[31\]\[25\] vssd1 vssd1 vccd1 vccd1 net2053
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06504__C net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09970_ net216 net2488 net418 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__mux2_1
Xhold748 total_design.core.regFile.register\[11\]\[13\] vssd1 vssd1 vccd1 vccd1 net2064
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06603__A2 _02092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold759 total_design.core.regFile.register\[2\]\[5\] vssd1 vssd1 vccd1 vccd1 net2075
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12137__B1 _05838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08921_ _04173_ _04174_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__and2_1
XANTENNA_wire458_X net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08852_ net968 _02029_ net533 vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__a21o_1
Xhold1404 total_design.core.regFile.register\[21\]\[13\] vssd1 vssd1 vccd1 vccd1 net2720
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06520__B net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1415 total_design.core.regFile.register\[27\]\[16\] vssd1 vssd1 vccd1 vccd1 net2731
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07803_ total_design.core.regFile.register\[1\]\[24\] net590 net571 total_design.core.regFile.register\[17\]\[24\]
+ _03305_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1426 total_design.core.regFile.register\[31\]\[31\] vssd1 vssd1 vccd1 vccd1 net2742
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1437 total_design.core.regFile.register\[21\]\[1\] vssd1 vssd1 vccd1 vccd1 net2753
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08783_ _02613_ net310 vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__nor2_1
Xhold1448 total_design.core.regFile.register\[21\]\[7\] vssd1 vssd1 vccd1 vccd1 net2764
+ sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_49_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1459 total_design.core.regFile.register\[6\]\[10\] vssd1 vssd1 vccd1 vccd1 net2775
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07734_ total_design.core.regFile.register\[28\]\[23\] net853 net763 total_design.core.regFile.register\[6\]\[23\]
+ _03241_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_140_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09323__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07665_ _03162_ _03165_ _03166_ _03175_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10469__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09550__C _04780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ _02940_ net504 net446 _02938_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_49_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06616_ _02182_ net462 vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__xor2_4
XTAP_TAPCELL_ROW_49_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07596_ total_design.core.regFile.register\[15\]\[20\] net604 _03109_ net686 vssd1
+ vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07619__A1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09335_ net321 _04386_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__nor2_1
X_06547_ total_design.core.regFile.register\[26\]\[1\] net925 net916 net913 vssd1
+ vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout140_X net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1261_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout617_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ net313 net298 _04296_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__or3_1
X_06478_ net744 net728 net727 vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08217_ net1352 net545 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[0\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_44_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09197_ net968 _02489_ _02490_ net537 vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_105_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08182__B _03375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09993__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ total_design.core.regFile.register\[2\]\[31\] net637 net609 total_design.core.regFile.register\[18\]\[31\]
+ _03627_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__a221o_1
XFILLER_0_161_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06414__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload180 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 clkload180/Y sky130_fd_sc_hd__clkinv_4
X_08079_ total_design.core.regFile.register\[9\]\[30\] net852 net800 total_design.core.regFile.register\[29\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12128__B1 _05826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10110_ net193 net2689 net402 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11090_ _01727_ _05030_ net350 net180 net520 vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_8_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ net202 net2203 net411 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold20 total_design.core.data_mem.data_read_adr_reg\[8\] vssd1 vssd1 vccd1 vccd1
+ net1336 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07555__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 total_design.core.data_mem.data_read_adr_reg\[24\] vssd1 vssd1 vccd1 vccd1
+ net1347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 total_design.core.math.pc_val\[3\] vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 total_design.core.data_mem.data_cpu_i_reg\[31\] vssd1 vssd1 vccd1 vccd1 net1369
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 total_design.core.data_mem.data_bus_i_reg\[9\] vssd1 vssd1 vccd1 vccd1 net1380
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold75 total_design.core.data_mem.data_cpu_i_reg\[18\] vssd1 vssd1 vccd1 vccd1 net1391
+ sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ clknet_leaf_75_clk total_design.core.data_mem.data_cpu_i\[9\] net1215 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[9\] sky130_fd_sc_hd__dfrtp_1
Xhold86 total_design.core.data_mem.data_cpu_i_reg\[19\] vssd1 vssd1 vccd1 vccd1 net1402
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 total_design.core.instr_mem.instruction_adr_stored\[18\] vssd1 vssd1 vccd1
+ vccd1 net1413 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11103__A1 total_design.core.data_bus_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11992_ total_design.lcd_display.row_2\[24\] _05832_ _05835_ total_design.lcd_display.row_2\[56\]
+ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__a22o_1
X_10943_ _05174_ _05201_ _05175_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__o21ai_1
X_13731_ clknet_leaf_75_clk total_design.core.data_mem.stored_write_data\[6\] net1220
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_97_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10379__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10874_ total_design.core.data_bus_o\[6\] net698 vssd1 vssd1 vccd1 vccd1 _05133_
+ sky130_fd_sc_hd__nand2_1
X_13662_ clknet_leaf_63_clk total_design.core.data_mem.data_read_adr_i\[2\] net1129
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06158__A total_design.core.ctrl.instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_156_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12613_ clknet_leaf_116_clk _00080_ net1212 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ clknet_leaf_37_clk total_design.core.data_mem.data_bus_i\[29\] net1070 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12544_ net1397 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12475_ net980 total_design.core.instr_mem.instruction_i\[1\] vssd1 vssd1 vccd1 vccd1
+ _01692_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14214_ clknet_leaf_78_clk _01394_ net1217 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfrtp_1
X_11426_ net1553 _05627_ net159 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__mux2_1
XANTENNA_6 _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14145_ clknet_leaf_42_clk _01325_ net1083 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11357_ _05355_ _05606_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12119__B1 _05848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10308_ net237 net2787 net494 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__mux2_1
X_14076_ clknet_leaf_109_clk _01256_ net1228 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[94\]
+ sky130_fd_sc_hd__dfrtp_1
X_11288_ _05509_ _05510_ _05512_ _05545_ _05546_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__08338__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13027_ clknet_leaf_16_clk _00494_ net1023 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10239_ net252 net2781 net502 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__mux2_1
XANTENNA__06340__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1040 net1045 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__buf_2
Xfanout1051 net1059 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__buf_2
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07010__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1062 net1065 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__clkbuf_2
Xfanout1073 net1074 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11673__S net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1084 net1105 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__buf_2
Xfanout1095 net1096 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13929_ clknet_leaf_94_clk _01109_ net1256 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10289__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07450_ total_design.core.regFile.register\[30\]\[17\] net838 net779 total_design.core.regFile.register\[27\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06401_ total_design.core.regFile.register\[29\]\[0\] net928 net947 _01950_ vssd1
+ vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__and4_1
XFILLER_0_123_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07381_ total_design.core.regFile.register\[13\]\[16\] net668 net564 total_design.core.regFile.register\[3\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a22o_1
X_09120_ _04353_ _04368_ _04369_ net450 vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10605__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06332_ wishbone.curr_state\[2\] wishbone.curr_state\[1\] vssd1 vssd1 vccd1 vccd1
+ _01911_ sky130_fd_sc_hd__nor2_2
XFILLER_0_127_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07077__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12070__A2 _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09471__B1 _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09051_ _04297_ _04302_ net316 vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__mux2_1
X_06263_ total_design.core.instr_mem.instruction_adr_i\[23\] total_design.core.instr_mem.instruction_adr_stored\[23\]
+ net981 vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__mux2_1
XANTENNA__06824__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08002_ total_design.core.regFile.register\[19\]\[28\] net641 net609 total_design.core.regFile.register\[18\]\[28\]
+ _03498_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold501 net51 vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
X_06194_ total_design.core.mem_ctrl.state\[1\] _01725_ total_design.core.mem_ctrl.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__and3b_1
XFILLER_0_13_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold512 total_design.lcd_display.row_2\[122\] vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold523 total_design.data_in_BUS\[30\] vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 net76 vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 total_design.core.mem_ctrl.next_next_fetch vssd1 vssd1 vccd1 vccd1 net1861
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold556 total_design.lcd_display.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08730__B net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07785__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 total_design.core.regFile.register\[31\]\[16\] vssd1 vssd1 vccd1 vccd1 net1883
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold578 total_design.core.regFile.register\[24\]\[0\] vssd1 vssd1 vccd1 vccd1 net1894
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 total_design.core.regFile.register\[27\]\[13\] vssd1 vssd1 vccd1 vccd1 net1905
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ net244 net2674 net418 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_115_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08904_ _02337_ _04099_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__nor2_1
X_09884_ net284 net2312 net426 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1107_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07537__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12530__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07914__X _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1201 total_design.core.regFile.register\[22\]\[9\] vssd1 vssd1 vccd1 vccd1 net2517
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 total_design.core.regFile.register\[20\]\[23\] vssd1 vssd1 vccd1 vccd1 net2528
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1223 total_design.core.regFile.register\[31\]\[3\] vssd1 vssd1 vccd1 vccd1 net2539
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ _04016_ _04018_ _04019_ _04021_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__o22a_1
Xhold1234 total_design.core.regFile.register\[14\]\[11\] vssd1 vssd1 vccd1 vccd1 net2550
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11583__S net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11436__X _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1245 total_design.core.regFile.register\[11\]\[2\] vssd1 vssd1 vccd1 vccd1 net2561
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout567_A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1256 total_design.core.regFile.register\[29\]\[10\] vssd1 vssd1 vccd1 vccd1 net2572
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 total_design.keypad0.counter\[6\] vssd1 vssd1 vccd1 vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ _03350_ _03369_ _04018_ _04020_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__a211o_1
Xhold1278 total_design.core.regFile.register\[24\]\[26\] vssd1 vssd1 vccd1 vccd1 net2594
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1289 total_design.core.regFile.register\[16\]\[28\] vssd1 vssd1 vccd1 vccd1 net2605
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07717_ total_design.core.regFile.register\[0\]\[22\] net684 _03222_ _03225_ vssd1
+ vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__o22a_4
XFILLER_0_135_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08697_ _03955_ net1925 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout355_X net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout734_A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08177__B _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09988__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07648_ total_design.core.regFile.register\[2\]\[21\] net637 _03158_ vssd1 vssd1
+ vccd1 vccd1 _03159_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06409__C net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout901_A _02016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ _03087_ _03089_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout1264_X net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09318_ _04548_ _04553_ _04559_ _04124_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_157_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12061__A2 _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ net167 net2051 net372 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09249_ total_design.core.math.pc_val\[9\] _04471_ vssd1 vssd1 vccd1 vccd1 _04494_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06815__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12260_ _06099_ _06100_ _06098_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_160_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ _05469_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12191_ _04399_ _06040_ net995 vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__mux2_1
XANTENNA__10662__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06579__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__clkbuf_4
X_11142_ _05400_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__inv_2
XANTENNA__07240__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__clkbuf_4
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA__06987__A_N _02515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__clkbuf_4
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
X_11073_ total_design.core.data_bus_o\[23\] total_design.core.data_bus_o\[31\] total_design.core.data_bus_o\[15\]
+ net699 net517 vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__a41o_1
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07528__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07824__X _03329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ net280 total_design.core.regFile.register\[21\]\[4\] net410 vssd1 vssd1 vccd1
+ vccd1 _00331_ sky130_fd_sc_hd__mux2_1
XANTENNA__11493__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08639__Y _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06751__A1 total_design.core.ctrl.instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_76_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11975_ net474 _05836_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__nor2_4
XFILLER_0_169_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09898__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13714_ clknet_leaf_27_clk total_design.core.data_mem.stored_read_data\[21\] net1077
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[21\] sky130_fd_sc_hd__dfrtp_1
X_10926_ net521 _05184_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07700__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13645_ clknet_leaf_49_clk total_design.core.data_mem.data_write_adr_i\[17\] net1101
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[17\] sky130_fd_sc_hd__dfrtp_1
X_10857_ _05096_ _05098_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07059__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10788_ net1266 total_design.core.data_bus_o\[7\] _05028_ vssd1 vssd1 vccd1 vccd1
+ _05047_ sky130_fd_sc_hd__and3_1
X_13576_ clknet_leaf_36_clk total_design.core.data_mem.data_bus_i\[12\] net1078 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[12\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09453__B1 _04290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06616__A _02182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12527_ net979 total_design.core.instr_mem.instruction_i\[27\] vssd1 vssd1 vccd1
+ vccd1 _01718_ sky130_fd_sc_hd__and2b_1
XFILLER_0_109_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12458_ net1904 net176 net345 vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__mux2_1
XANTENNA__11668__S net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11409_ _05663_ _05665_ _05667_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__and3_1
XANTENNA__10572__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12389_ total_design.core.math.pc_val\[27\] net988 vssd1 vssd1 vccd1 vccd1 _01649_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07767__B1 total_design.core.ctrl.imm_32\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07231__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14128_ clknet_leaf_109_clk _01308_ net1226 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_06950_ total_design.core.regFile.register\[10\]\[8\] net617 net579 total_design.core.regFile.register\[27\]\[8\]
+ _02498_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__a221o_1
X_14059_ clknet_leaf_91_clk _01239_ net1263 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12512__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06501__D net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06881_ total_design.core.regFile.register\[0\]\[6\] net876 _02423_ _02437_ vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[6\] sky130_fd_sc_hd__o22a_4
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08620_ total_design.lcd_display.cnt_20ms\[3\] _03910_ vssd1 vssd1 vccd1 vccd1 _03912_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ _03889_ _03893_ _03898_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__a21oi_1
X_07502_ total_design.core.regFile.register\[10\]\[18\] net837 net798 total_design.core.regFile.register\[29\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08482_ _03832_ _03833_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_46_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07298__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12291__A2 _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09692__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07433_ total_design.core.regFile.register\[1\]\[17\] net589 net585 total_design.core.regFile.register\[28\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08284__Y _03676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07364_ _02849_ _02892_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__xnor2_4
XANTENNA__12043__A2 _05810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09103_ net534 _04352_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__or2_1
XANTENNA__12247__B _02746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06315_ _01791_ _01798_ _01802_ _01849_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__or4b_1
XFILLER_0_165_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07295_ total_design.core.regFile.register\[19\]\[14\] net826 net801 total_design.core.regFile.register\[29\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09034_ net968 _02238_ _02239_ net537 vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_14_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1057_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06246_ net961 _01824_ _01823_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08741__A _03375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11578__S net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 total_design.lcd_display.row_1\[37\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10482__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06177_ net932 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__inv_2
Xhold331 total_design.lcd_display.row_2\[62\] vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06532__Y _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 total_design.lcd_display.row_1\[119\] vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07758__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1224_A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold353 net82 vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__C1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold364 total_design.lcd_display.row_2\[84\] vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold375 net78 vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06261__A _01771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07222__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold386 total_design.lcd_display.row_1\[65\] vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout684_A _02035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout800 net801 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__buf_4
Xhold397 total_design.lcd_display.row_2\[3\] vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 net813 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09936_ net216 net2558 net422 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__mux2_1
Xfanout822 _01966_ vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_8
Xfanout833 _01959_ vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__clkbuf_8
Xfanout844 net845 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_4
Xfanout855 _01947_ vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_8
Xfanout866 _01941_ vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__buf_2
XANTENNA__06411__D net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout877 net878 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__buf_2
X_09867_ net215 net2165 net430 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout851_A net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout888 _02023_ vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__buf_2
Xhold1020 total_design.core.regFile.register\[12\]\[23\] vssd1 vssd1 vccd1 vccd1 net2336
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout899 net900 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__buf_2
Xhold1031 total_design.core.regFile.register\[20\]\[16\] vssd1 vssd1 vccd1 vccd1 net2347
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 total_design.core.regFile.register\[17\]\[28\] vssd1 vssd1 vccd1 vccd1 net2358
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 total_design.core.regFile.register\[14\]\[24\] vssd1 vssd1 vccd1 vccd1 net2369
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ _04068_ _04070_ _04071_ _04072_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__or4b_1
X_09798_ net214 total_design.core.regFile.register\[28\]\[17\] net438 vssd1 vssd1
+ vccd1 vccd1 _00120_ sky130_fd_sc_hd__mux2_1
Xhold1064 total_design.core.regFile.register\[24\]\[5\] vssd1 vssd1 vccd1 vccd1 net2380
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1075 total_design.core.regFile.register\[29\]\[3\] vssd1 vssd1 vccd1 vccd1 net2391
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1086 total_design.core.regFile.register\[15\]\[10\] vssd1 vssd1 vccd1 vccd1 net2402
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06200__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1097 total_design.core.regFile.register\[10\]\[24\] vssd1 vssd1 vccd1 vccd1 net2413
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ _04003_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11760_ net516 _05693_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_159_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07289__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10711_ net209 net2250 net359 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11691_ net24 net937 _05690_ net2526 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__a22o_1
XANTENNA__10657__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout904_X net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13430_ clknet_leaf_156_clk _00897_ net1142 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10642_ net222 net2176 net478 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12034__A2 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13361_ clknet_leaf_151_clk _00828_ net1145 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10573_ net230 net2030 net370 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_172_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07997__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12312_ _01573_ _01575_ _06139_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07461__A2 _01932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13292_ clknet_leaf_174_clk _00759_ net1054 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11488__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12243_ _06082_ _06083_ _06085_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10392__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11545__A1 _05648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07749__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12174_ net902 _02292_ _06025_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06171__A total_design.core.data_cpu_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ _05379_ _05381_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__and2_1
X_11056_ net520 _05044_ _05054_ _05314_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__a31o_1
X_10007_ net202 net2842 net416 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11958_ _05802_ _05805_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__or2_4
XFILLER_0_80_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08826__A _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10909_ _05165_ _05167_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__nand2_1
XANTENNA__10567__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11889_ _05761_ _05765_ _05766_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__and3b_1
XFILLER_0_7_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06617__Y _02188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13628_ clknet_leaf_62_clk total_design.core.data_mem.data_write_adr_i\[0\] net1125
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12025__A2 _05832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13559_ clknet_leaf_164_clk _01026_ net1165 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11784__A1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07080_ _02619_ _02621_ _02623_ _02624_ vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__or4_2
XFILLER_0_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07452__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11536__A1 _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06512__C net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout129 net132 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_4
X_07982_ total_design.core.regFile.register\[15\]\[28\] net847 net777 total_design.core.regFile.register\[22\]\[28\]
+ _03479_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09721_ total_design.core.math.pc_val\[29\] _04905_ total_design.core.math.pc_val\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a21o_1
X_06933_ total_design.core.regFile.register\[0\]\[7\] net874 _02479_ _02486_ vssd1
+ vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__o22ai_1
X_09652_ net969 _03462_ _03464_ _04100_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__o211ai_1
X_06864_ total_design.core.regFile.register\[27\]\[6\] net781 net766 total_design.core.regFile.register\[6\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08603_ net2882 net338 net714 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[24\]
+ sky130_fd_sc_hd__and3_1
X_09583_ _03324_ net505 net448 _03323_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__o22a_1
XFILLER_0_171_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06795_ total_design.core.regFile.register\[31\]\[5\] net603 net595 total_design.core.regFile.register\[8\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08534_ total_design.data_in_BUS\[10\] net342 _03883_ vssd1 vssd1 vccd1 vccd1 _03884_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_26_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08465_ _03791_ _03794_ _03818_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__a21o_1
XANTENNA__10477__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout432_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1174_A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07416_ _02839_ _02843_ _02891_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__and3b_1
XFILLER_0_135_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08396_ total_design.keypad0.key_out\[6\] total_design.keypad0.key_out\[4\] _03715_
+ _03751_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12016__A2 _05804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07691__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07347_ total_design.core.regFile.register\[25\]\[15\] net844 _02875_ _02876_ vssd1
+ vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__a211o_1
XANTENNA__12421__C1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07979__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09567__A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07278_ _02805_ _02807_ _02809_ _02810_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout899_A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ net336 _03506_ _04269_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__o21bai_1
X_06229_ _01762_ _01772_ net1266 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__o21ai_4
XANTENNA__06651__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11527__A1 _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 total_design.core.data_mem.data_read_adr_reg2\[9\] vssd1 vssd1 vccd1 vccd1
+ net1466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 total_design.core.data_mem.data_read_adr_reg2\[20\] vssd1 vssd1 vccd1 vccd1
+ net1477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 total_design.core.data_mem.data_read_adr_reg2\[31\] vssd1 vssd1 vccd1 vccd1
+ net1488 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10225__B net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold183 total_design.core.math.pc_val\[19\] vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06422__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 total_design.core.data_mem.data_read_adr_reg2\[11\] vssd1 vssd1 vccd1 vccd1
+ net1510 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout630 net631 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_4
Xfanout641 net643 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_109_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09919_ net244 net1888 net425 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__mux2_1
Xfanout652 _02054_ vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout663 _02049_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_8
Xfanout674 net677 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout685 _02035_ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__buf_4
Xfanout696 net697 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_3_1_0_clk_X clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12930_ clknet_leaf_131_clk _00397_ net1197 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12861_ clknet_leaf_11_clk _00328_ net1020 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11812_ _05707_ net1874 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__nor2_1
X_12792_ clknet_leaf_135_clk _00259_ net1189 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10895__B net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14531_ net1303 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_68_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11743_ net1611 net959 net292 total_design.core.data_bus_o\[15\] vssd1 vssd1 vccd1
+ vccd1 _01371_ sky130_fd_sc_hd__a22o_1
XANTENNA__10387__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14462_ clknet_leaf_52_clk net1379 net1094 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12007__A2 _05804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11674_ _05609_ net1733 net130 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__mux2_1
XANTENNA__07682__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ clknet_leaf_115_clk _00880_ net1202 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10625_ _04119_ _04972_ _05002_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__or3_1
X_14393_ clknet_leaf_44_clk _01534_ vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_clk
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10556_ net170 net2821 net373 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__mux2_1
X_13344_ clknet_leaf_193_clk _00811_ net1013 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07434__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13275_ clknet_leaf_149_clk _00742_ net1149 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10487_ net183 net2017 net378 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__mux2_1
XANTENNA__11518__A1 _05651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12226_ _06068_ _06071_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12157_ net531 _05802_ _05813_ _05910_ _06010_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__o311a_1
XFILLER_0_102_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11108_ _01728_ _05030_ net515 total_design.core.data_bus_o\[12\] _05028_ vssd1 vssd1
+ vccd1 vccd1 _05367_ sky130_fd_sc_hd__o2111a_1
X_12088_ total_design.lcd_display.row_1\[116\] _05814_ _05829_ total_design.lcd_display.row_1\[108\]
+ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__a22o_1
XANTENNA__08147__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11039_ _05057_ _05297_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_34_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12494__A2 total_design.core.ctrl.instruction\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11681__S net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06580_ total_design.core.ctrl.instruction\[8\] _01918_ net888 net970 _02151_ vssd1
+ vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[1\] sky130_fd_sc_hd__a221o_2
XANTENNA__09647__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10297__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08250_ net1394 net557 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[0\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_60_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07201_ _02738_ _02718_ vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__nand2b_1
XANTENNA__06507__C net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08181_ net890 _03330_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[24\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11757__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07132_ total_design.core.regFile.register\[31\]\[11\] net831 _01986_ total_design.core.regFile.register\[2\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__a22o_1
XANTENNA__11757__B2 total_design.core.data_bus_o\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07063_ total_design.core.regFile.register\[28\]\[10\] net585 _02607_ net686 vssd1
+ vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__a211o_1
XANTENNA__11509__A1 _05609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12182__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10193__A0 _04401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ _03459_ _03460_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__or2_1
XANTENNA__08138__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ net506 _04928_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__and2_1
X_06916_ total_design.core.regFile.register\[14\]\[7\] net864 net845 total_design.core.regFile.register\[25\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__a22o_1
XANTENNA__09886__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07896_ total_design.core.regFile.register\[20\]\[26\] net671 net571 total_design.core.regFile.register\[17\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__a22o_1
XANTENNA__13322__RESET_B net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ _04861_ _04862_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__or2_1
XANTENNA__11693__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06847_ total_design.core.regFile.register\[25\]\[6\] net649 net587 total_design.core.regFile.register\[28\]\[6\]
+ _02403_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_104_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11591__S net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09638__B1 _04860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09566_ net296 _04434_ _04789_ _04796_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__o211a_1
X_06778_ _02335_ _02337_ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08517_ _03852_ _03867_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_121_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout814_A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ _04645_ _04730_ net326 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__mux2_1
XANTENNA__08185__B _03512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09996__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10000__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08448_ net931 _01759_ _03800_ _03801_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06417__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire305 _03642_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__buf_4
XFILLER_0_162_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08379_ total_design.keypad0.key_out\[3\] total_design.keypad0.key_out\[12\] vssd1
+ vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout602_X net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11748__B2 total_design.core.data_bus_o\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10410_ net224 net2228 net386 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11390_ _05643_ _05645_ _05646_ _05648_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06624__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10341_ net238 net2259 net490 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13060_ clknet_leaf_106_clk _00527_ net1233 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10272_ net249 net2548 net499 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12173__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12011_ total_design.lcd_display.row_2\[97\] _05846_ vssd1 vssd1 vccd1 vccd1 _05872_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11619__X _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10670__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09744__B _04966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout460 net461 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_2
Xfanout471 net473 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__buf_2
Xfanout482 _05011_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_8
X_13962_ clknet_leaf_86_clk _01142_ net1247 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout493 net494 vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11684__A0 _05630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09341__A2 _04581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ clknet_leaf_152_clk _00380_ net1146 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07203__A_N _02718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893_ clknet_leaf_85_clk _01073_ net1249 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11354__X _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12844_ clknet_leaf_165_clk _00311_ net1165 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12775_ clknet_leaf_173_clk _00242_ net1055 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08301__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14514_ net1286 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
X_11726_ _05692_ _01904_ net512 vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__and3b_1
XFILLER_0_12_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07655__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08852__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14445_ clknet_leaf_64_clk net1845 net1213 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06863__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11657_ _05624_ net1822 net131 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11739__B2 total_design.core.data_bus_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07407__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10608_ net224 net2074 net367 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__mux2_1
X_14376_ clknet_leaf_114_clk _01517_ net1204 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11588_ _05621_ net1701 net139 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__mux2_1
X_13327_ clknet_leaf_147_clk _00794_ net1152 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold908 total_design.core.regFile.register\[28\]\[11\] vssd1 vssd1 vccd1 vccd1 net2224
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold919 total_design.core.regFile.register\[0\]\[24\] vssd1 vssd1 vccd1 vccd1 net2235
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08080__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10539_ net238 net2189 net374 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06343__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13258_ clknet_leaf_25_clk _00725_ net1106 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12164__A1 net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11676__S net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12209_ net995 _04450_ net897 vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10580__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13189_ clknet_leaf_117_clk _00656_ net1161 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_07750_ total_design.core.regFile.register\[9\]\[23\] net663 net632 total_design.core.regFile.register\[16\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06701_ _02266_ vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[3\] sky130_fd_sc_hd__inv_2
XANTENNA__11675__A0 _05612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07681_ total_design.core.regFile.register\[12\]\[22\] net773 net771 total_design.core.regFile.register\[28\]\[22\]
+ _03190_ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06632_ total_design.core.regFile.register\[19\]\[2\] net824 net787 total_design.core.regFile.register\[13\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__a22o_1
X_09420_ net220 net2292 net455 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06358__X _01934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06563_ total_design.core.regFile.register\[15\]\[1\] net920 net911 net946 vssd1
+ vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__and4_1
X_09351_ _04590_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_950 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09096__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09096__B2 _01751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06518__B net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08302_ net1518 net940 _03685_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[8\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09282_ _02694_ net706 _04524_ _04105_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06494_ net743 net731 net723 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ net1433 net543 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[16\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_144_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout130_A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08733__B _02241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08164_ net893 _02492_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[7\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06534__A net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07115_ total_design.core.regFile.register\[21\]\[11\] net600 net592 total_design.core.regFile.register\[1\]\[11\]
+ _02656_ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__a221o_1
X_08095_ total_design.core.regFile.register\[5\]\[30\] net630 net579 total_design.core.regFile.register\[27\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08071__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload70 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA_fanout1137_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07046_ net966 net888 vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__nand2_1
Xclkload81 clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__inv_8
Xclkload92 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 clkload92/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_2_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout597_A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10490__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07365__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07031__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_145_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout764_A _01997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ net335 _03226_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__nor2_1
X_07948_ total_design.core.regFile.register\[25\]\[27\] net648 net629 total_design.core.regFile.register\[5\]\[27\]
+ _03444_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_3_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11666__A0 _05679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09580__A _04105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07879_ total_design.core.regFile.register\[15\]\[26\] net847 net824 total_design.core.regFile.register\[19\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09618_ _03418_ _04825_ _04844_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__or3_1
XFILLER_0_35_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06268__X _01847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ _05087_ _05123_ _05145_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__or3_1
XANTENNA__07885__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09549_ total_design.core.data_cpu_o\[22\] net754 vssd1 vssd1 vccd1 vccd1 _04781_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout817_X net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12560_ net1422 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12091__B1 _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07637__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08834__A1 total_design.core.data_mem.data_cpu_i\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11511_ net1520 _05628_ net151 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__mux2_1
XANTENNA__06845__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10665__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12491_ net979 total_design.core.instr_mem.instruction_i\[9\] vssd1 vssd1 vccd1 vccd1
+ _01700_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14230_ clknet_leaf_48_clk _01410_ net1103 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11442_ net1528 _05636_ net159 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__mux2_1
XANTENNA__06444__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11373_ _05049_ _05610_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__or2_2
XFILLER_0_1_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14161_ clknet_leaf_34_clk _01341_ net1066 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13112_ clknet_leaf_138_clk _00579_ net1185 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10324_ net175 net2344 net494 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__mux2_1
XANTENNA__07270__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14092_ clknet_leaf_99_clk _01272_ net1230 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11496__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13043_ clknet_leaf_178_clk _00510_ net1033 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10255_ net187 net2446 net501 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__mux2_1
XANTENNA__12181__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1200 net1201 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__clkbuf_4
Xfanout1211 net1212 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07022__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1222 net1265 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__buf_2
X_10186_ net161 total_design.core.regFile.register\[17\]\[31\] net395 vssd1 vssd1
+ vccd1 vccd1 _00486_ sky130_fd_sc_hd__mux2_1
Xfanout1233 net1235 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__clkbuf_4
Xfanout1244 net1246 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__clkbuf_4
Xfanout1255 net1256 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1266 net34 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__buf_4
Xfanout290 net291 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_2
XFILLER_0_89_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13945_ clknet_leaf_96_clk _01125_ net1254 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13876_ clknet_leaf_26_clk total_design.core.ctrl.imm_32\[15\] net1107 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[15\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07876__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12827_ clknet_leaf_143_clk _00294_ net1173 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12082__B1 _05826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07628__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12758_ clknet_leaf_153_clk _00225_ net1138 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11709_ net14 net934 net877 net2673 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__o22a_1
XANTENNA__10575__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12689_ clknet_leaf_148_clk _00156_ net1145 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14428_ clknet_leaf_32_clk total_design.core.data_out_INSTR\[23\] net1063 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06354__A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14359_ clknet_leaf_46_clk _00028_ net1088 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09250__A1 _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08053__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold705 total_design.core.regFile.register\[25\]\[19\] vssd1 vssd1 vccd1 vccd1 net2021
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09250__B2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold716 total_design.core.regFile.register\[27\]\[10\] vssd1 vssd1 vccd1 vccd1 net2032
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 total_design.core.regFile.register\[7\]\[23\] vssd1 vssd1 vccd1 vccd1 net2043
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold738 total_design.core.regFile.register\[9\]\[19\] vssd1 vssd1 vccd1 vccd1 net2054
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold749 total_design.core.regFile.register\[24\]\[11\] vssd1 vssd1 vccd1 vccd1 net2065
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07800__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08920_ net471 _03226_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07013__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ total_design.core.ctrl.instruction\[12\] total_design.core.ctrl.instruction\[14\]
+ _02029_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_51_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1405 total_design.core.regFile.register\[17\]\[24\] vssd1 vssd1 vccd1 vccd1 net2721
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 total_design.core.instr_mem.instruction_i\[6\] vssd1 vssd1 vccd1 vccd1 net2732
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07802_ total_design.core.regFile.register\[14\]\[24\] net625 net598 total_design.core.regFile.register\[21\]\[24\]
+ _03306_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__a221o_1
Xhold1427 total_design.core.regFile.register\[17\]\[7\] vssd1 vssd1 vccd1 vccd1 net2743
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1438 total_design.core.regFile.register\[23\]\[26\] vssd1 vssd1 vccd1 vccd1 net2754
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08782_ _02565_ total_design.core.data_mem.data_cpu_i\[9\] vssd1 vssd1 vccd1 vccd1
+ _04037_ sky130_fd_sc_hd__nor2_1
Xhold1449 total_design.core.regFile.register\[31\]\[7\] vssd1 vssd1 vccd1 vccd1 net2765
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11648__A0 _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07733_ total_design.core.regFile.register\[9\]\[23\] net850 net786 total_design.core.regFile.register\[13\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout178_A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ _03168_ _03170_ _03172_ _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__or4_1
X_09403_ _02944_ net701 _04640_ net533 vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__a211o_1
XFILLER_0_172_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06615_ _02185_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09069__A1 _02292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07595_ total_design.core.regFile.register\[11\]\[20\] net612 net585 total_design.core.regFile.register\[28\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__a22o_1
XANTENNA__08794__A_N total_design.core.data_mem.data_cpu_i\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06546_ total_design.core.regFile.register\[27\]\[1\] net925 net913 net911 vssd1
+ vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__and4_1
X_09334_ _04391_ _04574_ net319 vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07619__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09265_ _04193_ _04508_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__nand2_1
XANTENNA__10485__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06477_ total_design.core.regFile.register\[30\]\[0\] net747 net731 net727 vssd1
+ vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__and4_1
XFILLER_0_173_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08292__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13800__D total_design.core.data_mem.data_cpu_i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08216_ net561 net883 vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09196_ _04331_ _04442_ net327 vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__mux2_1
XANTENNA__06264__A _01771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12376__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08147_ total_design.core.regFile.register\[30\]\[31\] net660 net641 total_design.core.regFile.register\[19\]\[31\]
+ _03626_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__a221o_1
XANTENNA__08044__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload170 clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 clkload170/Y sky130_fd_sc_hd__bufinv_16
X_08078_ total_design.core.regFile.register\[12\]\[30\] net773 net771 total_design.core.regFile.register\[28\]\[30\]
+ _03571_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__a221o_1
Xclkload181 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 clkload181/Y sky130_fd_sc_hd__inv_8
XANTENNA_fanout881_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout979_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07029_ total_design.core.regFile.register\[18\]\[9\] net859 net814 total_design.core.regFile.register\[4\]\[9\]
+ net693 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_112_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ net205 net2792 net410 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__mux2_1
XANTENNA__07004__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06203__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold10 total_design.core.data_mem.data_read_adr_reg\[20\] vssd1 vssd1 vccd1 vccd1
+ net1326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 total_design.core.data_mem.data_read_adr_reg\[12\] vssd1 vssd1 vccd1 vccd1
+ net1337 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 total_design.core.data_mem.data_read_adr_reg\[30\] vssd1 vssd1 vccd1 vccd1
+ net1348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 total_design.core.data_mem.data_cpu_i_reg\[3\] vssd1 vssd1 vccd1 vccd1 net1359
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 total_design.core.data_mem.data_bus_i_reg\[6\] vssd1 vssd1 vccd1 vccd1 net1370
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 total_design.core.data_mem.data_cpu_i_reg\[27\] vssd1 vssd1 vccd1 vccd1 net1381
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__A0 _05652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold76 total_design.core.data_mem.data_cpu_i_reg\[20\] vssd1 vssd1 vccd1 vccd1 net1392
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold87 total_design.core.data_mem.data_bus_i_reg\[14\] vssd1 vssd1 vccd1 vccd1 net1403
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 total_design.core.instr_mem.instruction_adr_stored\[16\] vssd1 vssd1 vccd1
+ vccd1 net1414 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ net474 _05851_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__nor2_4
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13730_ clknet_leaf_74_clk total_design.core.data_mem.stored_write_data\[5\] net1220
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[5\] sky130_fd_sc_hd__dfrtp_2
X_10942_ _05165_ _05167_ _05171_ _05150_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__a31oi_1
XANTENNA__12637__RESET_B net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07858__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13661_ clknet_leaf_62_clk total_design.core.data_mem.data_read_adr_i\[1\] net1128
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[1\] sky130_fd_sc_hd__dfrtp_1
X_10873_ _05114_ _05117_ _05131_ _05112_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_78_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06530__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12612_ clknet_leaf_105_clk _00079_ net1233 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12064__B1 _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13592_ clknet_leaf_34_clk total_design.core.data_mem.data_bus_i\[28\] net1068 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06818__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12543_ net1410 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10395__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06294__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07491__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12474_ net982 total_design.core.ctrl.instruction\[0\] net883 _01691_ vssd1 vssd1
+ vccd1 vccd1 _01539_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213_ clknet_leaf_78_clk _01393_ net1217 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfrtp_1
X_11425_ net1583 _05677_ net157 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_7 _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14144_ clknet_leaf_43_clk _01324_ net1082 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07243__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11356_ _05606_ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10307_ net240 net2493 net495 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__mux2_1
X_14075_ clknet_leaf_91_clk _01255_ net1263 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[93\]
+ sky130_fd_sc_hd__dfrtp_1
X_11287_ _05488_ _05505_ _05541_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__and3_1
X_13026_ clknet_leaf_127_clk _00493_ net1191 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10238_ net263 net2668 net502 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__mux2_1
Xfanout1030 net1031 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07546__B2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1041 net1045 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__clkbuf_4
Xfanout1052 net1058 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__clkbuf_4
X_10169_ net232 net2071 net397 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1063 net1064 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__clkbuf_4
Xfanout1074 net1075 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__buf_2
Xfanout1085 net1105 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_4
Xfanout1096 net1105 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09299__A1 total_design.core.data_cpu_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09299__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13928_ clknet_leaf_83_clk _01108_ net1241 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07849__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_164_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13859_ clknet_leaf_47_clk total_design.core.mem_ctrl.next_state\[2\] net1089 vssd1
+ vssd1 vccd1 vccd1 total_design.core.mem_ctrl.state\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06400_ net926 net946 net909 vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__and3_1
XANTENNA__12055__B1 _05812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07380_ total_design.core.regFile.register\[10\]\[16\] net618 net575 total_design.core.regFile.register\[24\]\[16\]
+ _02906_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06331_ _01907_ _01909_ wishbone.curr_state\[0\] vssd1 vssd1 vccd1 vccd1 _01910_
+ sky130_fd_sc_hd__or3b_1
XANTENNA__06809__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_179_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08283__B net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09050_ _04300_ _04301_ net324 vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__mux2_1
X_06262_ total_design.core.data_adr_o\[17\] net962 vssd1 vssd1 vccd1 vccd1 _01841_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07482__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08001_ total_design.core.regFile.register\[20\]\[28\] net671 net571 total_design.core.regFile.register\[17\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__a22o_1
X_06193_ total_design.core.mem_ctrl.state\[2\] _01761_ vssd1 vssd1 vccd1 vccd1 _01773_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09223__A1 _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08026__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold502 total_design.keypad0.counter\[13\] vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold513 total_design.lcd_display.row_1\[50\] vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 net104 vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07234__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06371__X _01947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold535 total_design.lcd_display.row_2\[33\] vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 total_design.core.regFile.register\[20\]\[1\] vssd1 vssd1 vccd1 vccd1 net1862
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 total_design.lcd_display.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 total_design.core.regFile.register\[8\]\[1\] vssd1 vssd1 vccd1 vccd1 net1884
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 total_design.core.regFile.register\[31\]\[1\] vssd1 vssd1 vccd1 vccd1 net1895
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ net285 net2840 net418 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08903_ _04155_ _04156_ net312 _04142_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ _04115_ _04976_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout295_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 total_design.core.regFile.register\[28\]\[14\] vssd1 vssd1 vccd1 vccd1 net2518
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ total_design.core.data_mem.data_cpu_i\[30\] _03596_ _04025_ _04088_ _04024_
+ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__a311o_1
Xhold1213 total_design.core.regFile.register\[1\]\[6\] vssd1 vssd1 vccd1 vccd1 net2529
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10541__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08739__A _03090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1002_A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06745__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1224 total_design.core.regFile.register\[16\]\[25\] vssd1 vssd1 vccd1 vccd1 net2540
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 total_design.core.regFile.register\[30\]\[25\] vssd1 vssd1 vccd1 vccd1 net2551
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 total_design.core.regFile.register\[3\]\[15\] vssd1 vssd1 vccd1 vccd1 net2562
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 total_design.core.regFile.register\[20\]\[9\] vssd1 vssd1 vccd1 vccd1 net2573
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ _03395_ _03415_ _04016_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__a21bo_1
Xhold1268 total_design.core.regFile.register\[7\]\[16\] vssd1 vssd1 vccd1 vccd1 net2584
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout462_A _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06760__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1279 total_design.core.regFile.register\[7\]\[11\] vssd1 vssd1 vccd1 vccd1 net2595
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11165__A _05411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07716_ _03209_ _03213_ _03214_ _03224_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__or4_1
XANTENNA__07362__B _02868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08696_ total_design.keypad0.counter\[10\] _03954_ net1924 vssd1 vssd1 vccd1 vccd1
+ _03966_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07647_ total_design.core.regFile.register\[7\]\[21\] net653 net578 total_design.core.regFile.register\[27\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__a22o_1
XANTENNA__12046__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06409__D _01950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07578_ _03092_ vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[20\] sky130_fd_sc_hd__inv_2
XFILLER_0_82_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09317_ _04191_ _04554_ _04555_ _04558_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_118_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06529_ total_design.core.regFile.register\[16\]\[0\] net633 _02063_ _02086_ _02088_
+ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_91_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09462__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ _04481_ _04486_ _04492_ net451 vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__a31o_1
XFILLER_0_51_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08017__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09179_ net272 net2011 net456 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11210_ net302 _05461_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07225__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12190_ _06036_ _06039_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11141_ _05391_ _05395_ _05397_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_101_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__clkbuf_4
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__clkbuf_4
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__clkbuf_4
X_11072_ _05057_ _05221_ _05287_ _05288_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__a22o_1
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__clkbuf_4
X_10023_ net271 total_design.core.regFile.register\[21\]\[3\] net411 vssd1 vssd1 vccd1
+ vccd1 _00330_ sky130_fd_sc_hd__mux2_1
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11088__A1 total_design.core.data_bus_o\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08489__C1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11974_ _05799_ _05811_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__or2_2
X_13713_ clknet_leaf_27_clk total_design.core.data_mem.stored_read_data\[20\] net1073
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[20\] sky130_fd_sc_hd__dfrtp_1
X_10925_ total_design.core.data_bus_o\[4\] net698 vssd1 vssd1 vccd1 vccd1 _05184_
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_86_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13644_ clknet_leaf_56_clk total_design.core.data_mem.data_write_adr_i\[16\] net1113
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10856_ _05111_ _05112_ _05108_ _05109_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_27_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13575_ clknet_leaf_36_clk total_design.core.data_mem.data_bus_i\[11\] net1071 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[11\] sky130_fd_sc_hd__dfrtp_1
X_10787_ net520 net350 vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__nand2_1
XANTENNA__06175__Y _01757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09453__B2 _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12526_ net975 total_design.core.ctrl.instruction\[26\] net883 _01717_ vssd1 vssd1
+ vccd1 vccd1 _01565_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12457_ net2182 net183 net345 vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output91_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ net302 _05598_ _05653_ _05666_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__a31oi_4
XTAP_TAPCELL_ROW_10_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07216__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06191__X _01771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12388_ _01639_ _01644_ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__and2_1
XANTENNA__07767__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14127_ clknet_leaf_84_clk _01307_ net1245 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11339_ _05463_ _05597_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14058_ clknet_leaf_86_clk _01238_ net1248 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11684__S net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ clknet_leaf_152_clk _00476_ net1146 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06880_ _02429_ _02431_ _02433_ _02436_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__or4_1
XANTENNA__09154__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06742__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08550_ _03886_ _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__xor2_1
XANTENNA__08846__X _04101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07501_ total_design.core.regFile.register\[23\]\[18\] net810 net759 total_design.core.regFile.register\[21\]\[18\]
+ _03021_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__a221o_1
X_08481_ _03830_ _03831_ _03833_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_46_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07432_ total_design.core.regFile.register\[23\]\[17\] net678 net569 total_design.core.regFile.register\[17\]\[17\]
+ _02955_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07363_ _02890_ _02891_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_21_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09102_ _02342_ _04351_ net706 vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06314_ _01811_ _01814_ _01827_ _01892_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__and4_1
XANTENNA__07455__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07294_ total_design.core.regFile.register\[10\]\[14\] net837 _02825_ _02826_ vssd1
+ vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__a211o_1
XFILLER_0_150_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06245_ total_design.core.instr_mem.instruction_adr_i\[16\] total_design.core.instr_mem.instruction_adr_stored\[16\]
+ net985 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__mux2_1
X_09033_ _02241_ _04284_ net706 vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09396__Y _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08741__B _03421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold310 total_design.keypad0.counter\[0\] vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
X_06176_ total_design.keypad0.key_out\[13\] vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__inv_2
Xhold321 total_design.lcd_display.row_2\[35\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 net88 vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 total_design.lcd_display.row_2\[80\] vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold354 total_design.lcd_display.row_1\[47\] vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 total_design.lcd_display.row_1\[94\] vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold376 total_design.lcd_display.row_2\[90\] vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 total_design.lcd_display.row_2\[2\] vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout801 _01976_ vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__clkbuf_4
Xhold398 total_design.core.regFile.register\[15\]\[1\] vssd1 vssd1 vccd1 vccd1 net1714
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09935_ net213 total_design.core.regFile.register\[24\]\[17\] net422 vssd1 vssd1
+ vccd1 vccd1 _00248_ sky130_fd_sc_hd__mux2_1
Xfanout812 net813 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__buf_4
Xfanout823 net826 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout834 net837 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11594__S net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout845 _01954_ vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__buf_4
XANTENNA__06981__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout856 _01947_ vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__clkbuf_4
Xfanout867 _01941_ vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__clkbuf_8
X_09866_ net220 net2409 net432 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__mux2_1
Xfanout878 _05691_ vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__buf_2
Xhold1010 total_design.core.regFile.register\[3\]\[19\] vssd1 vssd1 vccd1 vccd1 net2326
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 total_design.core.regFile.register\[14\]\[12\] vssd1 vssd1 vccd1 vccd1 net2337
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 _02023_ vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09064__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1032 total_design.core.regFile.register\[4\]\[1\] vssd1 vssd1 vccd1 vccd1 net2348
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ _02468_ net458 vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__or2_1
Xhold1043 total_design.core.regFile.register\[1\]\[31\] vssd1 vssd1 vccd1 vccd1 net2359
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ net222 net2361 net440 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout844_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1054 total_design.core.regFile.register\[13\]\[15\] vssd1 vssd1 vccd1 vccd1 net2370
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08188__B _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06733__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1065 total_design.core.regFile.register\[6\]\[27\] vssd1 vssd1 vccd1 vccd1 net2381
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 total_design.core.regFile.register\[2\]\[23\] vssd1 vssd1 vccd1 vccd1 net2392
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09999__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10003__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1087 total_design.core.regFile.register\[5\]\[9\] vssd1 vssd1 vccd1 vccd1 net2403
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ _03112_ net457 total_design.core.data_mem.data_cpu_i\[21\] net299 vssd1 vssd1
+ vccd1 vccd1 _04003_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_107_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 total_design.core.regFile.register\[23\]\[19\] vssd1 vssd1 vccd1 vccd1 net2414
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08679_ total_design.keypad0.counter\[12\] _03955_ vssd1 vssd1 vccd1 vccd1 _03956_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_159_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09683__A1 _01757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout632_X net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12019__B1 _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10710_ net219 net2425 net357 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__mux2_1
XANTENNA__11490__A1 _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11690_ net13 net937 net879 net2202 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__a22o_1
X_10641_ net225 net2562 net478 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13360_ clknet_leaf_186_clk _00827_ net1038 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07446__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10572_ net238 net2193 net372 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_165_Right_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08932__A _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11793__A2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12311_ _01579_ total_design.core.math.pc_val\[18\] net522 vssd1 vssd1 vccd1 vccd1
+ _01488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10673__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13291_ clknet_leaf_115_clk _00758_ net1202 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12242_ _06083_ _06085_ _06082_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06452__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08946__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ net994 _04345_ _04346_ _06024_ net897 vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__o311a_1
XFILLER_0_31_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11124_ _05359_ _05371_ _05375_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__and3b_1
XFILLER_0_101_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06972__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11055_ _05243_ _05279_ _05294_ _05304_ net352 vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__o41a_1
XFILLER_0_155_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10006_ net207 net2003 net414 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09123__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11957_ _05799_ net474 _05813_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__nor3_4
XTAP_TAPCELL_ROW_28_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08826__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10908_ _05166_ _05143_ _05144_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__mux2_2
XANTENNA__11481__A1 _05645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11888_ _05765_ _05766_ _05761_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_117_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13627_ clknet_leaf_55_clk net1335 net1114 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10839_ _05085_ _05097_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_8__f_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_41_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07437__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13558_ clknet_leaf_160_clk _01025_ net1150 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06914__X _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08842__A total_design.core.ctrl.instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11679__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12509_ net975 total_design.core.instr_mem.instruction_i\[18\] vssd1 vssd1 vccd1
+ vccd1 _01709_ sky130_fd_sc_hd__and2b_1
XFILLER_0_140_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10583__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13489_ clknet_leaf_151_clk _00956_ net1146 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06362__A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06512__D net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07981_ total_design.core.regFile.register\[14\]\[28\] net862 net858 total_design.core.regFile.register\[18\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__a22o_1
XANTENNA__06963__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ total_design.core.math.pc_val\[29\] total_design.core.math.pc_val\[30\] _04905_
+ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__and3_1
X_06932_ _02481_ _02482_ _02483_ _02485_ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__or4_1
X_09651_ net322 _04877_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__or2_1
X_06863_ total_design.core.regFile.register\[20\]\[6\] net817 net812 total_design.core.regFile.register\[23\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08602_ total_design.data_in_BUS\[23\] net340 net715 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[23\]
+ sky130_fd_sc_hd__and3_1
X_09582_ _04768_ _04811_ net465 vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__mux2_1
X_06794_ total_design.core.regFile.register\[13\]\[5\] net668 net638 total_design.core.regFile.register\[2\]\[5\]
+ _02353_ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__a221o_1
XFILLER_0_171_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08533_ _03869_ _03871_ _03881_ _03882_ _03768_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_26_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout160_A _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__A2 _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09665__A1 _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08464_ _03816_ _03817_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_102_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07140__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07415_ _02939_ _02940_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__nor2_2
XFILLER_0_174_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08395_ total_design.keypad0.key_out\[5\] total_design.keypad0.key_out\[7\] vssd1
+ vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07428__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07346_ total_design.core.regFile.register\[14\]\[15\] net863 net835 total_design.core.regFile.register\[10\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08752__A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09200__X _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11589__S net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07277_ total_design.core.regFile.register\[19\]\[14\] net643 net627 total_design.core.regFile.register\[14\]\[14\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__a221o_1
XANTENNA__09567__B _04797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09016_ net472 _03459_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__nor2_1
X_06228_ _01762_ _01772_ net1266 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout794_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 total_design.core.data_mem.data_read_adr_reg2\[15\] vssd1 vssd1 vccd1 vccd1
+ net1456 sky130_fd_sc_hd__dlygate4sd3_1
X_06159_ total_design.core.ctrl.instruction\[16\] vssd1 vssd1 vccd1 vccd1 _01742_
+ sky130_fd_sc_hd__inv_2
Xhold151 total_design.core.data_mem.data_read_adr_reg2\[4\] vssd1 vssd1 vccd1 vccd1
+ net1467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 total_design.core.data_mem.state\[2\] vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold173 total_design.lcd_display.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 total_design.core.data_mem.data_read_adr_reg2\[24\] vssd1 vssd1 vccd1 vccd1
+ net1500 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07600__B1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06422__D net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold195 total_design.lcd_display.row_1\[20\] vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08943__A3 _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout961_A _01770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout582_X net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 net623 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__clkbuf_8
Xfanout631 _02062_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__buf_4
XANTENNA__06954__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout642 net643 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_4
X_09918_ net285 net1894 net425 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12488__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout653 _02054_ vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_109_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout664 net665 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__clkbuf_8
Xfanout675 net677 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__clkbuf_8
Xfanout686 net689 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06211__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout697 net700 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__buf_2
X_09849_ _04115_ _04974_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__nand2_1
XANTENNA__06706__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_X net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ clknet_4_1__leaf_clk _00327_ net1075 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07390__X _02917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11811_ total_design.lcd_display.cnt_20ms\[7\] _05705_ net1873 vssd1 vssd1 vccd1
+ vccd1 _05708_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12791_ clknet_leaf_123_clk _00258_ net1166 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10668__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ net1302 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
X_11742_ net1691 net957 net290 total_design.core.data_bus_o\[14\] vssd1 vssd1 vccd1
+ vccd1 _01370_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11463__A1 _05663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07131__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14437__Q total_design.core.instr_fetch vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14461_ clknet_leaf_52_clk net1452 net1094 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11673_ _05636_ net1747 net131 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13412_ clknet_leaf_106_clk _00879_ net1223 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10624_ net164 net2384 net366 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14392_ clknet_leaf_150_clk _01533_ net1148 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_133_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11499__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13343_ clknet_leaf_182_clk _00810_ net1040 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10555_ net173 net2739 net375 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__mux2_1
XANTENNA__08092__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13274_ clknet_leaf_133_clk _00741_ net1195 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ net185 net2460 net378 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12225_ _06069_ _06070_ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07565__X total_design.core.data_mem.data_cpu_i\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09592__B1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ _05823_ _05970_ _05994_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__nor3_1
X_11107_ total_design.core.data_bus_o\[11\] total_design.core.data_bus_o\[12\] total_design.core.data_bus_o\[13\]
+ net698 net511 vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__a41o_1
XFILLER_0_75_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12087_ _05938_ _05940_ _05942_ _05944_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_142_Left_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11038_ _05212_ _05237_ _05296_ _05215_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_34_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10578__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12989_ clknet_leaf_9_clk _00456_ net1019 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07658__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06357__A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07122__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_180_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_180_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_60_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Left_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07200_ net552 total_design.core.data_mem.data_cpu_i\[12\] total_design.core.ctrl.imm_32\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08180_ net890 _03282_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[23\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06644__X total_design.core.ctrl.imm_32\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11757__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07131_ total_design.core.regFile.register\[20\]\[11\] net818 net813 total_design.core.regFile.register\[23\]\[11\]
+ _02672_ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07062_ total_design.core.regFile.register\[9\]\[10\] net663 net597 total_design.core.regFile.register\[21\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__a22o_1
XANTENNA__07830__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07189__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4__f_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09583__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07475__X total_design.core.ctrl.imm_32\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_160_Left_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07964_ _03462_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09703_ total_design.core.data_cpu_o\[29\] net754 _04924_ _04927_ vssd1 vssd1 vccd1
+ vccd1 _04928_ sky130_fd_sc_hd__a211o_2
X_06915_ total_design.core.regFile.register\[11\]\[7\] net797 _01980_ total_design.core.regFile.register\[12\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__a22o_1
X_07895_ net553 _03395_ _03179_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11872__S net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_A _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ total_design.core.math.pc_val\[26\] _04838_ vssd1 vssd1 vccd1 vccd1 _04862_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07897__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06846_ total_design.core.regFile.register\[9\]\[6\] net665 net610 total_design.core.regFile.register\[18\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10488__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09565_ _04623_ _04687_ _04791_ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout542_A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09638__A1 total_design.core.data_cpu_o\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06777_ _02334_ _02338_ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__nand2_2
XANTENNA__13803__D total_design.core.data_mem.data_cpu_i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_136_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11445__A1 _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08516_ _03844_ _03864_ _03865_ _03866_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_121_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07649__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09496_ _04690_ _04729_ net461 vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__mux2_1
XANTENNA__07113__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11996__A2 _05812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08447_ _01758_ total_design.keypad0.key_out\[15\] vssd1 vssd1 vccd1 vccd1 _03801_
+ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_171_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_171_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout807_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09578__A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire306 _03551_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_4
X_08378_ total_design.keypad0.key_out\[3\] total_design.keypad0.key_out\[12\] vssd1
+ vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08074__B1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07329_ total_design.core.regFile.register\[20\]\[15\] net672 net579 total_design.core.regFile.register\[27\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__a22o_1
XANTENNA__06273__Y _01852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07098__A total_design.core.ctrl.instruction\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_143_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10340_ net241 net2100 net488 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout797_X net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10271_ net262 total_design.core.regFile.register\[14\]\[8\] net499 vssd1 vssd1 vccd1
+ vccd1 _00559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12010_ net2466 net709 _05862_ _05871_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06927__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout450 net451 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_4
Xfanout461 net462 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_2
Xfanout472 net473 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_2
X_13961_ clknet_leaf_93_clk _01141_ net1255 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout483 _05011_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_4
Xfanout494 net495 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__buf_6
X_12912_ clknet_leaf_186_clk _00379_ net1030 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07888__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13892_ clknet_leaf_110_clk _01072_ net1209 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09252__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07352__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12843_ clknet_leaf_120_clk _00310_ net1170 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10398__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_15__f_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774_ clknet_leaf_201_clk _00241_ net1004 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14513_ net1285 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_51_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13032__RESET_B net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11725_ net2854 net953 _05694_ vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_162_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_162_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08852__A2 _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14444_ clknet_leaf_64_clk net1631 net1213 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11656_ _05635_ net1713 net130 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10607_ net234 net2773 net368 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__mux2_1
X_14375_ clknet_leaf_20_clk _01516_ net1050 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11587_ _05477_ net1752 net137 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13326_ clknet_leaf_188_clk _00793_ net1028 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09000__B _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold909 total_design.core.regFile.register\[2\]\[20\] vssd1 vssd1 vccd1 vccd1 net2225
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07812__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10538_ net242 net2289 net373 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06343__C total_design.core.ctrl.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13257_ clknet_leaf_4_clk _00724_ net1033 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10469_ net263 total_design.core.regFile.register\[8\]\[8\] net379 vssd1 vssd1 vccd1
+ vccd1 _00751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12164__A2 _01766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12208_ _06053_ _06054_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_36_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13188_ clknet_leaf_105_clk _00655_ net1233 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06918__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _05754_ _05851_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_53_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07591__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06700_ net965 _02020_ _02265_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_84_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07680_ total_design.core.regFile.register\[17\]\[22\] net820 net814 total_design.core.regFile.register\[4\]\[22\]
+ net692 vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__a221o_1
XANTENNA__07879__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07343__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06631_ total_design.core.regFile.register\[31\]\[2\] net832 net760 total_design.core.regFile.register\[21\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11427__A1 _05663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09350_ _02770_ _02790_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06562_ total_design.core.regFile.register\[30\]\[1\] net925 net916 net946 vssd1
+ vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__and4_1
XANTENNA__10101__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08301_ total_design.core.data_mem.data_write_adr_reg\[8\] net548 net540 total_design.core.data_mem.data_read_adr_reg\[8\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__a221o_1
X_09281_ _02693_ _04522_ _04523_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_153_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_153_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06493_ total_design.core.regFile.register\[4\]\[0\] _02031_ net738 net734 vssd1
+ vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__and4_1
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08232_ net1868 net542 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[15\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_118_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06374__X _01950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08733__C _02292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08163_ net893 _02442_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07114_ total_design.core.regFile.register\[7\]\[11\] net652 net580 total_design.core.regFile.register\[27\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__a22o_1
XANTENNA__07803__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08094_ total_design.core.regFile.register\[30\]\[30\] net661 _03584_ _03585_ _03586_
+ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload60 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__clkinv_8
Xclkload71 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_77_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07045_ total_design.core.ctrl.instruction\[30\] _02028_ vssd1 vssd1 vccd1 vccd1
+ _02591_ sky130_fd_sc_hd__nand2_1
Xclkload82 clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 clkload82/Y sky130_fd_sc_hd__inv_8
XFILLER_0_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1032_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload93 clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_149_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12155__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07646__A _03157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06909__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout492_A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07365__B _02893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ _04247_ _04248_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_145_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07582__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07947_ total_design.core.regFile.register\[11\]\[27\] net614 net567 total_design.core.regFile.register\[12\]\[27\]
+ _03445_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_3_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06790__B1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07878_ total_design.core.regFile.register\[30\]\[26\] net839 _03378_ _03379_ vssd1
+ vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__a211o_1
XANTENNA__07334__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ _04825_ _04844_ _03418_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06829_ _02388_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[5\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_74_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11418__A1 _05477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ net904 _04779_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__or2_1
XANTENNA__10011__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09800__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09479_ _04704_ _04713_ net449 vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_144_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_144_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ net1589 _05612_ net149 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12490_ net980 total_design.core.ctrl.instruction\[8\] net882 _01699_ vssd1 vssd1
+ vccd1 vccd1 _01547_ sky130_fd_sc_hd__a22o_1
XANTENNA__06725__A _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11441_ net1523 _05652_ net160 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08047__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09795__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14160_ clknet_leaf_34_clk _01340_ net1066 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11372_ _05358_ _05628_ _05629_ _05630_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__and4b_1
XFILLER_0_132_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13111_ clknet_leaf_162_clk _00578_ net1166 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10323_ net176 net2050 net493 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__mux2_1
X_14091_ clknet_leaf_89_clk _01271_ net1261 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10681__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12146__A2 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ clknet_leaf_146_clk _00509_ net1178 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10254_ net189 net2434 net501 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1201 net1265 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__buf_2
Xfanout1212 net1265 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10185_ net165 net1964 net396 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1223 net1224 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__clkbuf_4
Xfanout1234 net1235 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__buf_2
Xfanout1245 net1246 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__clkbuf_4
Xfanout1256 net1257 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout280 net283 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_2
Xfanout291 net292 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__dlymetal6s2s_1
X_13944_ clknet_leaf_74_clk _01124_ net1220 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07325__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13875_ clknet_leaf_26_clk total_design.core.ctrl.imm_32\[14\] net1107 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06619__B net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12826_ clknet_leaf_125_clk _00293_ net1188 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07089__A1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12757_ clknet_leaf_156_clk _00224_ net1142 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_135_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_135_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11708_ net12 net936 net879 net2870 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12688_ clknet_leaf_189_clk _00155_ net1030 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08038__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14427_ clknet_leaf_29_clk total_design.core.data_out_INSTR\[22\] net1063 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[22\] sky130_fd_sc_hd__dfrtp_1
X_11639_ _05652_ net1646 net134 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14358_ clknet_leaf_46_clk _00027_ net1088 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09250__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11593__A0 _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold706 total_design.core.regFile.register\[25\]\[31\] vssd1 vssd1 vccd1 vccd1 net2022
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold717 total_design.core.regFile.register\[20\]\[27\] vssd1 vssd1 vccd1 vccd1 net2033
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold728 total_design.core.regFile.register\[30\]\[4\] vssd1 vssd1 vccd1 vccd1 net2044
+ sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ clknet_leaf_11_clk _00776_ net1025 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10591__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold739 total_design.core.regFile.register\[10\]\[28\] vssd1 vssd1 vccd1 vccd1 net2055
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ clknet_leaf_109_clk _01465_ net1228 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06641__Y _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12137__A2 _05812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08850_ total_design.core.ctrl.instruction\[12\] total_design.core.ctrl.instruction\[14\]
+ _02029_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_51_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07801_ total_design.core.regFile.register\[5\]\[24\] net629 net586 total_design.core.regFile.register\[28\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__a22o_1
XANTENNA__07564__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1406 total_design.core.regFile.register\[31\]\[8\] vssd1 vssd1 vccd1 vccd1 net2722
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08761__A1 _03395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08761__B2 _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1417 total_design.core.regFile.register\[4\]\[4\] vssd1 vssd1 vccd1 vccd1 net2733
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08781_ total_design.core.data_mem.data_cpu_i\[13\] _02770_ vssd1 vssd1 vccd1 vccd1
+ _04036_ sky130_fd_sc_hd__and2b_1
Xhold1428 total_design.core.regFile.register\[11\]\[14\] vssd1 vssd1 vccd1 vccd1 net2744
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1439 total_design.core.regFile.register\[28\]\[30\] vssd1 vssd1 vccd1 vccd1 net2755
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07732_ total_design.core.regFile.register\[31\]\[23\] net831 net794 total_design.core.regFile.register\[11\]\[23\]
+ _03239_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_140_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07663_ total_design.core.regFile.register\[8\]\[21\] net594 _03173_ net687 vssd1
+ vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__a211o_1
XANTENNA__13704__Q total_design.core.data_cpu_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09402_ _04638_ _04639_ net706 vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06614_ net461 _02182_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__and2b_1
XANTENNA__09069__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07594_ _03101_ _03103_ _03105_ _03107_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__or4_1
X_09333_ _04483_ _04573_ net331 vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__mux2_1
X_06545_ net752 _02118_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[0\]
+ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_126_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout338_A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09264_ _04289_ _04506_ net317 vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06476_ net744 net730 net726 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06545__A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08215_ total_design.core.data_mem.state\[1\] total_design.core.data_mem.state\[2\]
+ _01749_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__and3b_1
XFILLER_0_117_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08029__B1 _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09195_ _04441_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1247_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12376__A2 _03375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ total_design.core.regFile.register\[28\]\[31\] net586 _03636_ net687 vssd1
+ vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11584__A0 _05651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11597__S net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload160 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 clkload160/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_31_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08077_ total_design.core.regFile.register\[20\]\[30\] net816 net814 total_design.core.regFile.register\[4\]\[30\]
+ net693 vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__a221o_1
Xclkload171 clknet_leaf_84_clk vssd1 vssd1 vccd1 vccd1 clkload171/Y sky130_fd_sc_hd__clkinv_2
Xclkload182 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 clkload182/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__12128__A2 _05812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07028_ total_design.core.regFile.register\[21\]\[9\] net761 _02573_ _02575_ vssd1
+ vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__a211o_1
XANTENNA__06280__A net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_A _01934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10006__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold11 total_design.core.data_mem.data_read_adr_reg\[17\] vssd1 vssd1 vccd1 vccd1
+ net1327 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07555__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 total_design.core.data_mem.data_read_adr_reg\[4\] vssd1 vssd1 vccd1 vccd1
+ net1338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 total_design.core.data_mem.data_read_adr_reg\[3\] vssd1 vssd1 vccd1 vccd1
+ net1349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 total_design.core.math.pc_val\[11\] vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08979_ net334 _02234_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__nor2_1
XANTENNA__06763__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 total_design.core.data_mem.data_cpu_i_reg\[17\] vssd1 vssd1 vccd1 vccd1 net1371
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08919__B _03273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold66 total_design.core.mem_ctrl.state\[0\] vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 total_design.core.data_mem.data_bus_i_reg\[10\] vssd1 vssd1 vccd1 vccd1 net1393
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _05755_ _05851_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__nor2_4
Xhold88 total_design.core.math.pc_val\[16\] vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 total_design.bus_full vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11103__A3 _05049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12300__A2 _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ _05195_ _05196_ _05198_ _05180_ _05177_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__a2111o_1
X_13660_ clknet_leaf_62_clk total_design.core.data_mem.data_read_adr_i\[0\] net1128
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10872_ _05115_ _05117_ _05111_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ clknet_leaf_6_clk _00078_ net1017 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ clknet_leaf_34_clk total_design.core.data_mem.data_bus_i\[27\] net1068 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[27\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10676__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_117_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12542_ net1399 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06294__A2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12473_ net982 total_design.core.instr_mem.instruction_i\[0\] vssd1 vssd1 vccd1 vccd1
+ _01691_ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14212_ clknet_leaf_78_clk _01392_ net1217 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12367__A2 _03330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ _05358_ net302 _05625_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_50_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11575__A0 _05609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_8 _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ clknet_leaf_35_clk _01323_ net1068 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11355_ _05602_ _05471_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06461__Y _02035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12119__A2 _05840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07794__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ net253 total_design.core.regFile.register\[13\]\[10\] net492 vssd1 vssd1
+ vccd1 vccd1 _00593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14074_ clknet_leaf_87_clk _01254_ net1250 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06190__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11286_ _05540_ _05541_ _05505_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_67_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13025_ clknet_leaf_118_clk _00492_ net1169 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10237_ net267 net1886 net500 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__mux2_1
XANTENNA__08743__A1 _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1020 net1021 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07573__X _03090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1031 net1036 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09705__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1042 net1045 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__buf_2
X_10168_ net230 net2502 net397 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__mux2_1
Xfanout1053 net1054 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06754__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1064 net1065 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__buf_2
XFILLER_0_83_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1075 net1081 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__buf_2
Xfanout1086 net1105 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__buf_2
Xfanout1097 net1099 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09299__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10099_ net238 net2395 net403 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13927_ clknet_leaf_83_clk _01107_ net1243 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13858_ clknet_leaf_46_clk total_design.core.mem_ctrl.next_state\[1\] net1087 vssd1
+ vssd1 vccd1 vccd1 total_design.core.mem_ctrl.state\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_wire306_A _03551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10586__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12809_ clknet_leaf_14_clk _00276_ net1026 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_108_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13789_ clknet_leaf_59_clk total_design.core.data_mem.next_read net1127 vssd1 vssd1
+ vccd1 vccd1 total_design.core.data_mem.data_read sky130_fd_sc_hd__dfrtp_1
X_06330_ net1266 _01905_ _01908_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09471__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06261_ _01771_ _01839_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08000_ total_design.core.regFile.register\[15\]\[28\] net605 net583 total_design.core.regFile.register\[6\]\[28\]
+ _03496_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_96_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11566__A0 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06192_ net998 net997 total_design.core.instr_fetch vssd1 vssd1 vccd1 vccd1 _01772_
+ sky130_fd_sc_hd__or3_2
XFILLER_0_128_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold503 total_design.keypad0.counter\[10\] vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold514 total_design.lcd_display.row_2\[83\] vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold525 total_design.lcd_display.row_2\[27\] vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 total_design.data_in_BUS\[0\] vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 total_design.lcd_display.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07785__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ _04116_ _04972_ _04980_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__or3_1
Xhold558 _05708_ vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 total_design.core.regFile.register\[2\]\[1\] vssd1 vssd1 vccd1 vccd1 net1885
+ sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap288 _03092_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08902_ net324 _04149_ net316 vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _04968_ _04971_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09615__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07537__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12530__A2 total_design.core.ctrl.instruction\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08833_ _04029_ _04087_ _04026_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__o21a_1
Xhold1203 total_design.core.regFile.register\[25\]\[26\] vssd1 vssd1 vccd1 vccd1 net2519
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 total_design.core.regFile.register\[30\]\[22\] vssd1 vssd1 vccd1 vccd1 net2530
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 total_design.core.regFile.register\[13\]\[7\] vssd1 vssd1 vccd1 vccd1 net2541
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08739__B _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1236 total_design.core.regFile.register\[1\]\[23\] vssd1 vssd1 vccd1 vccd1 net2552
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 total_design.core.regFile.register\[17\]\[10\] vssd1 vssd1 vccd1 vccd1 net2563
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ net307 _03322_ _03350_ _03369_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__o22a_1
Xhold1258 total_design.core.regFile.register\[6\]\[17\] vssd1 vssd1 vccd1 vccd1 net2574
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 total_design.core.regFile.register\[17\]\[1\] vssd1 vssd1 vccd1 vccd1 net2585
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07715_ total_design.core.regFile.register\[7\]\[22\] net653 _03223_ net687 vssd1
+ vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__a211o_1
X_08695_ _03956_ _03965_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout455_A _04117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07646_ _03157_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[21\]
+ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07170__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10496__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07577_ _01748_ net885 net550 _03041_ total_design.core.ctrl.imm_32\[21\] vssd1 vssd1
+ vccd1 vccd1 _03092_ sky130_fd_sc_hd__o41ai_2
XANTENNA_fanout622_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ net313 net298 _04354_ _04557_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_24_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06528_ total_design.core.regFile.register\[7\]\[0\] net652 _02065_ _02073_ net689
+ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_63_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14265__Q total_design.core.math.pc_val\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09247_ net298 _04489_ _04490_ _04491_ _04488_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06459_ _01923_ net896 _02019_ _01744_ _01743_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09178_ _04121_ _04425_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__nor2_1
XANTENNA__11557__A0 _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08129_ _03609_ _03615_ _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__or3_2
XANTENNA__07818__B _03322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11140_ _05391_ _05395_ _05398_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__a21o_1
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10780__A1 total_design.core.data_bus_o\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__clkbuf_4
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09592__Y _04822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__clkbuf_4
X_11071_ net351 _05281_ _05290_ _05329_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__a31o_1
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07528__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ net278 net2511 net411 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__mux2_1
XANTENNA__06736__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06883__A_N net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ net531 _05799_ _05813_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__nor3_2
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10924_ _05153_ _05181_ _05182_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__a21bo_1
X_13712_ clknet_leaf_27_clk total_design.core.data_mem.stored_read_data\[19\] net1076
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[19\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07161__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07700__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13643_ clknet_leaf_58_clk total_design.core.data_mem.data_write_adr_i\[15\] net1118
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10855_ _05113_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13574_ clknet_leaf_38_clk total_design.core.data_mem.data_bus_i\[10\] net1078 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10786_ net517 net352 vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__nor2_2
XFILLER_0_137_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09453__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12525_ net975 total_design.core.instr_mem.instruction_i\[26\] vssd1 vssd1 vccd1
+ vccd1 _01717_ sky130_fd_sc_hd__and2b_1
XFILLER_0_125_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12456_ net2053 net185 net345 vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ _05360_ net304 vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12387_ total_design.core.math.pc_val\[26\] net523 _01646_ _01647_ vssd1 vssd1 vccd1
+ vccd1 _01496_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14126_ clknet_leaf_101_clk _01306_ net1236 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08964__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output84_A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11338_ _05530_ _05536_ _05590_ _05535_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14057_ clknet_leaf_97_clk _01237_ net1246 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[75\]
+ sky130_fd_sc_hd__dfrtp_1
X_11269_ _05524_ _05527_ _05525_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13008_ clknet_leaf_186_clk _00475_ net1031 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12512__A2 total_design.core.ctrl.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_158_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07500_ total_design.core.regFile.register\[26\]\[18\] net869 net819 total_design.core.regFile.register\[17\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__a22o_1
X_08480_ _03807_ _03811_ _03805_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_46_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07431_ total_design.core.regFile.register\[5\]\[17\] net628 net593 total_design.core.regFile.register\[8\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__a22o_1
XANTENNA_wire309_X net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07362_ _02889_ _02868_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_21_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ _02341_ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06313_ _01838_ _01847_ net929 _01836_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__and4b_1
XFILLER_0_162_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07293_ total_design.core.regFile.register\[11\]\[14\] net797 net762 total_design.core.regFile.register\[21\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09032_ _02240_ _04283_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__xnor2_1
X_06244_ total_design.core.data_mem.data_read total_design.core.data_mem.data_write
+ total_design.core.data_adr_o\[16\] vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08741__C _03512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold300 total_design.lcd_display.row_2\[63\] vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold311 total_design.lcd_display.row_1\[125\] vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
X_06175_ total_design.core.data_cpu_o\[28\] vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold322 total_design.lcd_display.row_2\[58\] vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10211__A0 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold333 total_design.lcd_display.row_2\[120\] vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07758__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08955__A1 _02188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold344 total_design.lcd_display.row_1\[14\] vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 total_design.lcd_display.row_2\[118\] vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 net102 vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06966__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 net42 vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11875__S net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold388 total_design.lcd_display.row_2\[45\] vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net805 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__clkbuf_8
Xhold399 total_design.lcd_display.row_2\[117\] vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ net221 net2269 net424 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1112_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout813 _01970_ vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__buf_4
Xfanout824 net826 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_37_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout835 net836 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__buf_4
Xfanout846 net849 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_8
Xfanout857 net860 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_8
X_09865_ net227 net2441 net432 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__mux2_1
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14517__1289 vssd1 vssd1 vccd1 vccd1 net1289 _14517__1289/LO sky130_fd_sc_hd__conb_1
XANTENNA__06718__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1000 total_design.core.regFile.register\[3\]\[25\] vssd1 vssd1 vccd1 vccd1 net2316
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08102__X _03595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout868 _01941_ vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__buf_4
XANTENNA_fanout572_A _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout879 _05690_ vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__buf_2
XANTENNA__13806__D total_design.core.data_mem.data_cpu_i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1011 total_design.core.regFile.register\[27\]\[11\] vssd1 vssd1 vccd1 vccd1 net2327
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1022 total_design.core.regFile.register\[8\]\[15\] vssd1 vssd1 vccd1 vccd1 net2338
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 total_design.core.regFile.register\[30\]\[14\] vssd1 vssd1 vccd1 vccd1 net2349
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ _02263_ _02286_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__nor2_1
Xhold1044 total_design.core.regFile.register\[2\]\[27\] vssd1 vssd1 vccd1 vccd1 net2360
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ net227 net1998 net440 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1055 total_design.core.regFile.register\[17\]\[15\] vssd1 vssd1 vccd1 vccd1 net2371
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 total_design.core.regFile.register\[17\]\[26\] vssd1 vssd1 vccd1 vccd1 net2382
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1077 total_design.core.regFile.register\[30\]\[27\] vssd1 vssd1 vccd1 vccd1 net2393
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ _02918_ total_design.core.data_mem.data_cpu_i\[16\] _02968_ net309 vssd1
+ vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__o2bb2a_1
Xhold1088 total_design.core.regFile.register\[14\]\[2\] vssd1 vssd1 vccd1 vccd1 net2404
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 total_design.core.regFile.register\[14\]\[18\] vssd1 vssd1 vccd1 vccd1 net2415
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09132__A1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ total_design.keypad0.counter\[10\] total_design.keypad0.counter\[11\] _03954_
+ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09683__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07629_ total_design.core.regFile.register\[12\]\[21\] net773 net771 total_design.core.regFile.register\[28\]\[21\]
+ _03140_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__a221o_1
XANTENNA__06276__Y _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_46_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10640_ net232 net2728 net479 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10571_ net240 net2607 net370 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__mux2_1
XANTENNA__08932__B _04101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12310_ net899 _03040_ _01578_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07997__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13290_ clknet_leaf_19_clk _00757_ net1049 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout994_X net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10526__Y _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12241_ total_design.core.math.pc_val\[11\] total_design.core.program_count.imm_val_reg\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06452__B _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08946__A1 total_design.core.math.pc_val\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07749__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_163_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ _06022_ _06023_ net994 vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__or3b_1
XFILLER_0_102_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11123_ _05359_ _05378_ _05375_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_55_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11054_ total_design.core.data_bus_o\[29\] net695 net352 _05305_ net518 vssd1 vssd1
+ vccd1 vccd1 _05313_ sky130_fd_sc_hd__a221o_1
XANTENNA__06709__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_178_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11702__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ net211 net2525 net416 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07382__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09123__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11373__X _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_101_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09123__B2 _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ net474 _05817_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_28_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07134__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10907_ _05127_ _05143_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__nand2_1
X_11887_ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10838_ _05076_ _05081_ _05083_ _05084_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__o211ai_1
X_13626_ clknet_leaf_55_clk net1348 net1114 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09003__B _02968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11769__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10769_ total_design.core.mem_ctrl.state\[1\] _01760_ vssd1 vssd1 vccd1 vccd1 _05028_
+ sky130_fd_sc_hd__nor2_4
XFILLER_0_137_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13557_ clknet_leaf_166_clk _01024_ net1157 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08842__B _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07988__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12508_ net974 total_design.core.ctrl.instruction\[17\] net881 _01708_ vssd1 vssd1
+ vccd1 vccd1 _01556_ sky130_fd_sc_hd__a22o_1
X_13488_ clknet_leaf_186_clk _00955_ net1036 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12439_ net2722 net262 net346 vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06660__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06362__B net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06948__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14109_ clknet_leaf_88_clk _01289_ net1249 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07745__Y _03253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07980_ total_design.core.regFile.register\[1\]\[28\] net829 net795 total_design.core.regFile.register\[11\]\[28\]
+ _03477_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09165__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06931_ total_design.core.regFile.register\[8\]\[7\] net805 _02484_ net691 vssd1
+ vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09650_ _04828_ _04875_ net468 vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__mux2_1
XANTENNA__10104__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06862_ total_design.core.regFile.register\[30\]\[6\] net840 net796 total_design.core.regFile.register\[11\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__a22o_1
XANTENNA__07373__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08601_ total_design.data_in_BUS\[22\] net340 net715 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[22\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__07912__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09581_ net471 _03322_ _04173_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__o21ai_1
X_06793_ total_design.core.regFile.register\[7\]\[5\] net654 net645 total_design.core.regFile.register\[26\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__a22o_1
XANTENNA__11724__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08532_ _03869_ _03871_ _03881_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07921__B _03421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07125__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08736__C _02746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ _03787_ _03815_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout153_A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07414_ _02917_ _02937_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_102_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08394_ total_design.data_in_BUS\[4\] _01888_ net519 vssd1 vssd1 vccd1 vccd1 _03750_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07345_ total_design.core.regFile.register\[16\]\[15\] net856 net778 total_design.core.regFile.register\[22\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout418_A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08752__B total_design.core.data_mem.data_cpu_i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07979__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07276_ total_design.core.regFile.register\[13\]\[14\] net669 net565 total_design.core.regFile.register\[3\]\[14\]
+ _02808_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09015_ _04267_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__inv_2
X_06227_ _01796_ _01780_ _01785_ _01805_ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__and4b_1
XFILLER_0_27_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06651__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold130 total_design.core.math.pc_val\[25\] vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09050__A0 _04300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold141 total_design.core.data_mem.data_bus_i_reg\[11\] vssd1 vssd1 vccd1 vccd1 net1457
+ sky130_fd_sc_hd__dlygate4sd3_1
X_06158_ total_design.core.ctrl.instruction\[15\] vssd1 vssd1 vccd1 vccd1 _01741_
+ sky130_fd_sc_hd__inv_2
Xhold152 total_design.core.instr_mem.instruction_adr_stored\[8\] vssd1 vssd1 vccd1
+ vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 total_design.core.data_mem.data_read_adr_reg2\[10\] vssd1 vssd1 vccd1 vccd1
+ net1479 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout787_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 total_design.core.data_mem.data_read_adr_reg2\[19\] vssd1 vssd1 vccd1 vccd1
+ net1490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold185 total_design.core.data_mem.data_read_adr_reg2\[30\] vssd1 vssd1 vccd1 vccd1
+ net1501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 total_design.lcd_display.row_1\[26\] vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 net611 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__clkbuf_4
Xfanout621 net622 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__buf_4
Xfanout632 _02061_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_8
X_09917_ _04115_ _04978_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__nand2_1
Xfanout643 _02058_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout954_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout575_X net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout654 _02054_ vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_97_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout665 _02049_ vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout676 net677 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10014__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout687 net689 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__buf_4
X_09848_ _04112_ _04971_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__nor2_1
Xfanout698 net699 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09803__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ net161 net2638 net444 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11810_ total_design.lcd_display.cnt_20ms\[7\] total_design.lcd_display.cnt_20ms\[8\]
+ _05705_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__and3_1
X_12790_ clknet_leaf_153_clk _00257_ net1138 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06728__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07116__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08313__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11999__B1 _05850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11741_ net1821 net956 _05059_ _05695_ vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06447__B _01915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11672_ _05652_ net1725 net130 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__mux2_1
X_14460_ clknet_leaf_39_clk net1592 net1091 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10623_ net165 net1919 net367 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__mux2_1
X_13411_ clknet_leaf_9_clk _00878_ net1020 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10684__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14391_ clknet_leaf_134_clk _01532_ net1190 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13342_ clknet_leaf_181_clk _00809_ net1043 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10554_ net177 net2381 net375 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__mux2_1
XANTENNA__14453__Q total_design.core.instr_mem.instruction_adr_i\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ clknet_leaf_195_clk _00740_ net1010 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10485_ net191 net2397 net378 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12224_ total_design.core.math.pc_val\[9\] total_design.core.program_count.imm_val_reg\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12155_ net2406 net710 _05999_ _06009_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11106_ _05363_ _05364_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__nor2_1
X_12086_ total_design.lcd_display.row_2\[76\] _05806_ _05812_ total_design.lcd_display.row_1\[92\]
+ _05943_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_88_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08147__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11037_ _05231_ _05233_ _05239_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_34_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07355__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12483__A_N net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07107__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12100__B1 _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12988_ clknet_leaf_12_clk _00455_ net1025 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_82_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11939_ _05754_ _05800_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06357__B _01932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13609_ clknet_leaf_58_clk net1330 net1117 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10594__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06881__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14516__1288 vssd1 vssd1 vccd1 vccd1 net1288 _14516__1288/LO sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_12_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07130_ total_design.core.regFile.register\[19\]\[11\] net826 net762 total_design.core.regFile.register\[21\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09280__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06373__A total_design.core.ctrl.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07061_ total_design.core.regFile.register\[22\]\[10\] net674 net593 total_design.core.regFile.register\[8\]\[10\]
+ _02605_ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09684__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07916__B _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ _03459_ _03460_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_79_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13707__Q total_design.core.data_cpu_o\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08138__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06914_ total_design.core.regFile.register\[0\]\[7\] net683 _02462_ _02467_ vssd1
+ vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__o22a_4
X_09702_ total_design.core.ctrl.instruction\[29\] net888 _04926_ net906 vssd1 vssd1
+ vccd1 vccd1 _04927_ sky130_fd_sc_hd__a22o_1
X_07894_ _03395_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[26\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__07346__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09633_ total_design.core.math.pc_val\[26\] _04838_ vssd1 vssd1 vccd1 vccd1 _04861_
+ sky130_fd_sc_hd__and2_1
X_06845_ total_design.core.regFile.register\[7\]\[6\] net654 net635 total_design.core.regFile.register\[16\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a22o_1
XANTENNA__11693__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09564_ _04195_ _04794_ _04664_ _04443_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__o2bb2a_1
X_06776_ _02108_ total_design.core.data_mem.data_cpu_i\[4\] _02336_ vssd1 vssd1 vccd1
+ vccd1 _02338_ sky130_fd_sc_hd__o21a_4
XANTENNA__09638__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08515_ _03850_ _03864_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_121_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09495_ net336 _03064_ _04176_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_121_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout156_X net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout535_A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08310__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08446_ _01758_ total_design.keypad0.key_out\[15\] vssd1 vssd1 vccd1 vccd1 _03800_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_93_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_173_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08377_ _03710_ _03734_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[2\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06872__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout702_A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire307 _03302_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06609__C1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07328_ total_design.core.regFile.register\[11\]\[15\] net614 net584 total_design.core.regFile.register\[6\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__a22o_1
XANTENNA__07806__D1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09271__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06624__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07098__B total_design.core.ctrl.instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07259_ _02791_ _02792_ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__nor2_1
XANTENNA__10009__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10270_ net267 net2262 net496 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07826__B _03330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07585__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08845__A_N total_design.core.ctrl.instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06222__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout440 net441 vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__clkbuf_8
Xfanout451 _04125_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_2
Xfanout462 _02184_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_4
X_13960_ clknet_leaf_82_clk _01140_ net1221 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[42\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout473 _02111_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_2
Xfanout484 _05007_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout495 _05005_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_4
X_12911_ clknet_leaf_160_clk _00378_ net1150 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10679__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13891_ clknet_leaf_88_clk _01071_ net1250 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[101\]
+ sky130_fd_sc_hd__dfrtp_1
X_12842_ clknet_leaf_21_clk _00309_ net1106 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12773_ clknet_leaf_119_clk _00240_ net1169 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08301__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14512_ net1284 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
X_11724_ net1 net953 vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__nor2_2
XFILLER_0_139_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14443_ clknet_leaf_77_clk net1728 net1216 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11655_ _05618_ net1703 net129 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__mux2_1
XANTENNA__06863__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10606_ net229 net2658 net368 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__mux2_1
X_11586_ _05478_ _05479_ _05674_ _05675_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__or4b_4
X_14374_ clknet_leaf_18_clk _01515_ net1051 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10537_ net255 net2775 net373 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__mux2_1
X_13325_ clknet_leaf_6_clk _00792_ net1017 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12149__B1 _05848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07576__X total_design.core.ctrl.imm_32\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10468_ _04452_ net2436 net377 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__mux2_1
XANTENNA__06480__X _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13256_ clknet_leaf_117_clk _00723_ net1162 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _06053_ _06054_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_36_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13187_ clknet_leaf_9_clk _00654_ net1016 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_max_cap333_A _02233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10399_ net282 net1967 net385 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__mux2_1
X_12138_ total_design.lcd_display.row_2\[79\] _05806_ _05815_ total_design.lcd_display.row_1\[87\]
+ _05992_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_53_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12069_ total_design.lcd_display.row_2\[51\] _05849_ _05852_ total_design.lcd_display.row_2\[11\]
+ _05927_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_1_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08848__A _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07328__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08200__X _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10589__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06630_ total_design.core.regFile.register\[9\]\[2\] net851 net806 total_design.core.regFile.register\[5\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__a22o_1
XANTENNA__07471__B _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06561_ total_design.core.regFile.register\[18\]\[1\] net925 net948 net916 vssd1
+ vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__and4_1
XFILLER_0_75_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08300_ net1472 net941 _03684_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[7\]
+ sky130_fd_sc_hd__o21a_1
X_09280_ _02693_ _04522_ net702 vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__a21oi_1
X_06492_ net742 net738 net734 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__and3_1
XANTENNA__07500__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08231_ net1403 net542 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[14\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__11721__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08162_ net893 _02395_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08870__X _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07113_ total_design.core.regFile.register\[5\]\[11\] net631 net601 total_design.core.regFile.register\[31\]\[11\]
+ _02650_ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12606__Q total_design.core.regFile.register\[29\]\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08093_ total_design.core.regFile.register\[25\]\[30\] net649 net595 total_design.core.regFile.register\[8\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__a22o_1
XANTENNA__06606__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload50 clknet_leaf_175_clk vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_70_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07044_ total_design.core.ctrl.instruction\[30\] _02541_ vssd1 vssd1 vccd1 vccd1
+ _02590_ sky130_fd_sc_hd__xor2_1
Xclkload61 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_77_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload72 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 clkload72/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__06831__A _02367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload83 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload94 clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 clkload94/Y sky130_fd_sc_hd__inv_12
XFILLER_0_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07567__B1 total_design.core.ctrl.imm_32\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06550__B net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1025_A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07031__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ net335 _03322_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_10_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout485_A _05007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07946_ total_design.core.regFile.register\[22\]\[27\] net676 net668 total_design.core.regFile.register\[13\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__a22o_1
XANTENNA__08758__A _03206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07877_ total_design.core.regFile.register\[24\]\[26\] net791 net787 total_design.core.regFile.register\[13\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__a22o_1
XANTENNA__10499__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout652_A _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ _03370_ _03369_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__and2b_1
X_06828_ total_design.core.regFile.register\[0\]\[5\] net876 _02372_ _02387_ vssd1
+ vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_168_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09547_ _04777_ _04778_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__or2_1
X_06759_ total_design.core.regFile.register\[27\]\[4\] net577 net573 total_design.core.regFile.register\[24\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10626__A0 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12091__A2 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ net295 _04327_ _04530_ _04687_ _04712_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08429_ _03780_ _03781_ _03779_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06845__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11440_ net1594 _05613_ net158 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__mux2_1
Xclkload0 clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_62_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06444__C _01915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11371_ total_design.core.data_bus_o\[31\] net699 net510 vssd1 vssd1 vccd1 vccd1
+ _05630_ sky130_fd_sc_hd__a21o_2
XFILLER_0_132_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09528__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13110_ clknet_leaf_154_clk _00577_ net1136 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10322_ net184 net2670 net493 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__mux2_1
X_14090_ clknet_leaf_86_clk _01270_ net1248 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07270__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13041_ clknet_leaf_160_clk _00508_ net1150 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10253_ net193 net2097 net500 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__mux2_1
XANTENNA__07558__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07022__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ net170 net2748 net394 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__mux2_1
Xfanout1202 net1204 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__clkbuf_4
Xfanout1213 net1214 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06230__A0 total_design.core.instr_mem.instruction_adr_i\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1224 net1240 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__clkbuf_4
Xfanout1235 net1240 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08939__Y _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1246 net1252 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1257 net1264 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__clkbuf_2
Xfanout270 net271 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515__1287 vssd1 vssd1 vccd1 vccd1 net1287 _14515__1287/LO sky130_fd_sc_hd__conb_1
Xfanout281 net283 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_2
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_2
X_13943_ clknet_leaf_82_clk _01123_ net1220 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10202__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13874_ clknet_leaf_68_clk total_design.core.ctrl.imm_32\[13\] net1109 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07730__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14178__Q net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ clknet_leaf_196_clk _00292_ net1009 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07089__A2 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12082__A2 _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12756_ clknet_leaf_141_clk _00223_ net1182 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06475__X _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11707_ net11 net936 net879 net1946 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__a22o_1
X_12687_ clknet_leaf_162_clk _00154_ net1153 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09011__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14426_ clknet_leaf_27_clk total_design.core.data_out_INSTR\[21\] net1076 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09235__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11638_ _05613_ net1651 net133 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14357_ clknet_leaf_45_clk _00026_ net1088 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11569_ _05680_ net1624 net143 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold707 total_design.core.regFile.register\[18\]\[3\] vssd1 vssd1 vccd1 vccd1 net2023
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold718 total_design.core.regFile.register\[28\]\[1\] vssd1 vssd1 vccd1 vccd1 net2034
+ sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ clknet_leaf_28_clk _00775_ net1074 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold729 total_design.core.regFile.register\[4\]\[21\] vssd1 vssd1 vccd1 vccd1 net2045
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14288_ clknet_leaf_98_clk _01464_ net1244 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13239_ clknet_leaf_162_clk _00706_ net1166 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07549__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07013__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07800_ total_design.core.regFile.register\[30\]\[24\] net660 net653 total_design.core.regFile.register\[7\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__a22o_1
XANTENNA__08761__A2 _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1407 total_design.core.regFile.register\[23\]\[8\] vssd1 vssd1 vccd1 vccd1 net2723
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08780_ _02818_ total_design.core.data_mem.data_cpu_i\[14\] vssd1 vssd1 vccd1 vccd1
+ _04035_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1418 total_design.core.regFile.register\[9\]\[8\] vssd1 vssd1 vccd1 vccd1 net2734
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1429 total_design.core.regFile.register\[26\]\[13\] vssd1 vssd1 vccd1 vccd1 net2745
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07731_ total_design.core.regFile.register\[19\]\[23\] net823 net802 total_design.core.regFile.register\[8\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07662_ total_design.core.regFile.register\[25\]\[21\] net648 net629 total_design.core.regFile.register\[5\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__a22o_1
XANTENNA__10112__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09901__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09401_ _02941_ _04617_ _04637_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__and3_1
X_06613_ net552 total_design.core.data_mem.data_cpu_i\[1\] total_design.core.ctrl.imm_32\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a21oi_4
X_07593_ total_design.core.regFile.register\[19\]\[20\] net640 net624 total_design.core.regFile.register\[14\]\[20\]
+ _03106_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06544_ _02112_ _02114_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__nor2_2
X_09332_ _04526_ _04572_ net463 vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__mux2_1
XANTENNA__12073__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09263_ _04506_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__inv_2
X_06475_ net741 net729 net724 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__and3_4
XANTENNA__13720__Q total_design.core.data_cpu_o\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06545__B _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08214_ _03658_ net561 _03657_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.next_write
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_62_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09194_ net463 _04440_ _04438_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08145_ total_design.core.regFile.register\[23\]\[31\] net679 net667 total_design.core.regFile.register\[13\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout400_A _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1142_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07788__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload150 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 clkload150/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_30_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08076_ total_design.core.regFile.register\[5\]\[30\] net808 _03566_ _03567_ _03569_
+ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__a2111o_1
Xclkload161 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 clkload161/Y sky130_fd_sc_hd__clkinv_4
Xclkload172 clknet_leaf_85_clk vssd1 vssd1 vccd1 vccd1 clkload172/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__13809__D total_design.core.data_mem.data_cpu_i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkload183 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 clkload183/Y sky130_fd_sc_hd__clkinv_2
X_07027_ total_design.core.regFile.register\[16\]\[9\] net856 net788 total_design.core.regFile.register\[13\]\[9\]
+ _02574_ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_8_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07004__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout867_A _01941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_X net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 total_design.core.data_mem.data_read_adr_reg\[6\] vssd1 vssd1 vccd1 vccd1
+ net1328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 total_design.core.data_mem.data_read_adr_reg\[27\] vssd1 vssd1 vccd1 vccd1
+ net1339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 total_design.core.data_mem.data_read_adr_reg\[16\] vssd1 vssd1 vccd1 vccd1
+ net1350 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10811__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08978_ _04224_ _04230_ net328 vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__mux2_1
Xhold45 total_design.core.data_mem.data_bus_i_reg\[5\] vssd1 vssd1 vccd1 vccd1 net1361
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 total_design.core.data_mem.data_cpu_i_reg\[2\] vssd1 vssd1 vccd1 vccd1 net1372
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 total_design.core.math.pc_val\[31\] vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ total_design.core.regFile.register\[19\]\[27\] net825 net800 total_design.core.regFile.register\[29\]\[27\]
+ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__a221o_1
Xhold78 total_design.core.data_mem.data_cpu_i_reg\[0\] vssd1 vssd1 vccd1 vccd1 net1394
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 total_design.core.data_mem.data_bus_i_reg\[13\] vssd1 vssd1 vccd1 vccd1 net1405
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10940_ _05177_ _05198_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__nor2_1
XANTENNA__10022__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07712__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09811__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10871_ _05111_ _05118_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12610_ clknet_leaf_131_clk _00077_ net1199 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12064__A2 _05830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13590_ clknet_leaf_34_clk total_design.core.data_mem.data_bus_i\[26\] net1067 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12541_ net1430 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06818__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_6__f_clk_X clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12472_ _01733_ _01690_ _01689_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_151_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07491__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14211_ clknet_leaf_60_clk _01391_ net1132 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11423_ net1630 _05626_ net159 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__mux2_1
XANTENNA__10692__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07779__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_9 _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14142_ clknet_leaf_43_clk _01322_ net1082 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11354_ _05457_ _05571_ _05608_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__or3b_4
XFILLER_0_85_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07243__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08015__X _03512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10305_ net251 net2198 net494 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__mux2_1
X_11285_ _05540_ _05541_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__nand2_1
X_14073_ clknet_leaf_96_clk _01253_ net1255 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06190__B net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12524__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13024_ clknet_leaf_193_clk _00491_ net1013 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10236_ net272 net2150 net502 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1010 net1015 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_4
Xfanout1021 net1027 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08743__A2 _03467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1032 net1036 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_4
X_10167_ net236 net2841 net396 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__mux2_1
Xfanout1043 net1045 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_4
Xfanout1054 net1058 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07951__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1065 net1081 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_156_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1076 net1080 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__clkbuf_4
Xfanout1087 net1089 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10098_ net242 net2241 net405 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1098 net1099 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__clkbuf_4
X_13926_ clknet_leaf_95_clk _01106_ net1254 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07703__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13857_ clknet_leaf_46_clk total_design.core.mem_ctrl.next_state\[0\] net1097 vssd1
+ vssd1 vccd1 vccd1 total_design.core.mem_ctrl.state\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12808_ clknet_leaf_23_clk _00275_ net1055 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12055__A2 _05810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13788_ clknet_leaf_56_clk total_design.core.data_mem.stored_data_adr\[31\] net1114
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[31\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08564__C net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06809__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12739_ clknet_leaf_5_clk _00206_ net1022 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06365__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06260_ total_design.core.instr_mem.instruction_adr_i\[17\] total_design.core.instr_mem.instruction_adr_stored\[17\]
+ net981 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07482__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08861__A total_design.core.instr_fetch vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14293__RESET_B net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14409_ clknet_leaf_41_clk total_design.core.data_out_INSTR\[4\] net1090 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06191_ net998 net997 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__or2_2
XFILLER_0_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold504 total_design.lcd_display.row_2\[106\] vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold515 total_design.lcd_display.row_2\[0\] vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold526 total_design.data_in_BUS\[4\] vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold537 total_design.core.regFile.register\[13\]\[1\] vssd1 vssd1 vccd1 vccd1 net1853
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold548 net96 vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold559 total_design.core.regFile.register\[31\]\[30\] vssd1 vssd1 vccd1 vccd1 net1875
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ total_design.core.ctrl.instruction\[10\] net556 total_design.core.ctrl.instruction\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__nand3b_2
XANTENNA__10107__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08901_ net459 _04152_ _04154_ net325 vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ net163 net2089 net431 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11727__A net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__C1 _04628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08832_ total_design.core.data_mem.data_cpu_i\[29\] net306 _04028_ vssd1 vssd1 vccd1
+ vccd1 _04087_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_57_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1204 total_design.core.regFile.register\[19\]\[9\] vssd1 vssd1 vccd1 vccd1 net2520
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1215 total_design.core.regFile.register\[21\]\[27\] vssd1 vssd1 vccd1 vccd1 net2531
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07942__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1226 total_design.core.regFile.register\[1\]\[26\] vssd1 vssd1 vccd1 vccd1 net2542
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08739__C _03187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1237 total_design.core.regFile.register\[18\]\[19\] vssd1 vssd1 vccd1 vccd1 net2553
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 total_design.core.regFile.register\[5\]\[0\] vssd1 vssd1 vccd1 vccd1 net2564
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ _03440_ _03459_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__and2_1
XFILLER_0_174_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout183_A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1259 total_design.core.regFile.register\[29\]\[6\] vssd1 vssd1 vccd1 vccd1 net2575
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09144__C1 _04101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07714_ total_design.core.regFile.register\[5\]\[22\] net629 net625 total_design.core.regFile.register\[14\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08694_ net2649 _03955_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07645_ total_design.core.regFile.register\[0\]\[21\] net875 _03144_ _03156_ vssd1
+ vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_68_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout448_A _04189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09203__Y _04450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12046__A2 _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07576_ total_design.core.ctrl.instruction\[31\] net885 _02149_ _03091_ net550 vssd1
+ vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[21\] sky130_fd_sc_hd__a221o_4
X_06527_ _02097_ _02098_ _02099_ _02100_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__or4_2
X_09315_ _02743_ net508 net446 _02739_ _04556_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__o221a_1
XFILLER_0_146_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ _02588_ _04102_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__nand2_1
X_06458_ _01923_ net896 _02019_ _01742_ _01741_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14514__1286 vssd1 vssd1 vccd1 vccd1 net1286 _14514__1286/LO sky130_fd_sc_hd__conb_1
X_09177_ _01753_ net752 _04424_ net905 _04423_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__o221a_4
X_06389_ total_design.core.regFile.register\[19\]\[0\] net927 net949 net912 vssd1
+ vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08128_ total_design.core.regFile.register\[13\]\[31\] net787 _03603_ _03618_ _03619_
+ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07225__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout984_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08059_ net306 _03552_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__or2_1
XANTENNA__10017__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10780__A2 total_design.core.data_bus_o\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__clkbuf_4
X_11070_ net520 _05291_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__nand2_1
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ net245 net2753 net410 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__mux2_1
XANTENNA__07933__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06230__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11972_ net474 _05833_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__nor2_4
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13711_ clknet_leaf_33_clk total_design.core.data_mem.stored_read_data\[18\] net1070
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[18\] sky130_fd_sc_hd__dfrtp_1
X_10923_ _05153_ _05155_ _05159_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__or3_1
XANTENNA__10687__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13642_ clknet_leaf_55_clk total_design.core.data_mem.data_write_adr_i\[14\] net1117
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[14\] sky130_fd_sc_hd__dfrtp_1
X_10854_ _05111_ _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__nor2_1
XANTENNA__12037__A2 _05838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13573_ clknet_leaf_35_clk total_design.core.data_mem.data_bus_i\[9\] net1071 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10785_ total_design.core.data_bus_o\[18\] net696 _05042_ net517 vssd1 vssd1 vccd1
+ vccd1 _05044_ sky130_fd_sc_hd__a211o_1
XFILLER_0_52_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12524_ net975 total_design.core.ctrl.instruction\[25\] net882 _01716_ vssd1 vssd1
+ vccd1 vccd1 _01564_ sky130_fd_sc_hd__a22o_1
XANTENNA__07464__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12455_ net2554 net189 net345 vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11548__A1 _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11406_ net302 _05594_ _05653_ _05664_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__a31oi_4
XTAP_TAPCELL_ROW_10_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07216__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12386_ net899 _03421_ net523 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_10_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14125_ clknet_leaf_88_clk _01305_ net1251 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11337_ _05595_ net294 _05537_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__or3b_2
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14056_ clknet_leaf_110_clk _01236_ net1225 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[74\]
+ sky130_fd_sc_hd__dfrtp_1
X_11268_ _05520_ _05526_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__and2_1
X_13007_ clknet_leaf_147_clk _00474_ net1150 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10219_ _04866_ net2657 net391 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11199_ _05042_ _05457_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07924__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08559__C net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13909_ clknet_leaf_92_clk _01089_ net1262 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10597__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07430_ total_design.core.regFile.register\[9\]\[17\] net663 net632 total_design.core.regFile.register\[16\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12028__A2 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07361_ _02868_ _02889_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__and2b_1
XFILLER_0_57_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06312_ _01817_ _01833_ _01889_ _01890_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__and4_1
XFILLER_0_150_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09100_ _02291_ _04317_ _04349_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_21_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07455__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07292_ total_design.core.regFile.register\[18\]\[14\] net857 net786 total_design.core.regFile.register\[13\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_135_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09031_ _02115_ _02187_ _04282_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__a21oi_2
X_06243_ _01808_ _01821_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11539__A1 _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06174_ total_design.core.data_cpu_o\[9\] vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold301 total_design.lcd_display.row_1\[25\] vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 total_design.lcd_display.row_2\[25\] vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 total_design.lcd_display.row_2\[68\] vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 total_design.lcd_display.row_2\[59\] vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08955__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 total_design.lcd_display.row_1\[36\] vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold356 total_design.lcd_display.row_2\[114\] vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 _01363_ vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 total_design.lcd_display.row_2\[123\] vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold389 total_design.lcd_display.row_2\[38\] vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ net225 net2629 net424 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout803 net805 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout814 net815 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__buf_4
Xfanout825 net826 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout398_A _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout836 net837 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout847 net849 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_8
X_09864_ net232 net2635 net433 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__mux2_1
Xfanout858 net859 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1105_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1001 total_design.core.regFile.register\[4\]\[26\] vssd1 vssd1 vccd1 vccd1 net2317
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout869 net872 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__clkbuf_8
Xhold1012 total_design.core.regFile.register\[9\]\[21\] vssd1 vssd1 vccd1 vccd1 net2328
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ total_design.core.data_mem.data_cpu_i\[0\] _02106_ _04069_ vssd1 vssd1 vccd1
+ vccd1 _04070_ sky130_fd_sc_hd__a21bo_1
Xhold1023 total_design.core.regFile.register\[15\]\[16\] vssd1 vssd1 vccd1 vccd1 net2339
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 total_design.core.regFile.register\[7\]\[21\] vssd1 vssd1 vccd1 vccd1 net2350
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ net234 net2518 net441 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1045 total_design.core.regFile.register\[28\]\[16\] vssd1 vssd1 vccd1 vccd1 net2361
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09117__C1 _04100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1056 total_design.core.regFile.register\[10\]\[6\] vssd1 vssd1 vccd1 vccd1 net2372
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 total_design.core.regFile.register\[16\]\[9\] vssd1 vssd1 vccd1 vccd1 net2383
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08746_ _03157_ _03178_ _03206_ _03226_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__o22a_1
Xhold1078 total_design.core.regFile.register\[13\]\[14\] vssd1 vssd1 vccd1 vccd1 net2394
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 total_design.core.regFile.register\[3\]\[12\] vssd1 vssd1 vccd1 vccd1 net2405
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07670__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ total_design.keypad0.counter\[8\] total_design.keypad0.counter\[9\] _03953_
+ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12019__A2 _05848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07628_ total_design.core.regFile.register\[30\]\[21\] net839 net814 total_design.core.regFile.register\[4\]\[21\]
+ net692 vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__a221o_1
XANTENNA__10300__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06351__C1 _01915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07559_ total_design.core.regFile.register\[17\]\[19\] net820 net803 total_design.core.regFile.register\[8\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ net253 net2782 net369 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07446__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06654__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09229_ net452 _04474_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12240_ total_design.core.math.pc_val\[11\] total_design.core.program_count.imm_val_reg\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06225__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12171_ _06020_ _06021_ _06012_ _06015_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__o211a_1
XANTENNA__08946__A2 _02014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11122_ _05380_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__inv_2
Xhold890 total_design.core.regFile.register\[9\]\[1\] vssd1 vssd1 vccd1 vccd1 net2206
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11053_ _05037_ _05046_ _05305_ net352 vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07906__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ net216 total_design.core.regFile.register\[22\]\[18\] net414 vssd1 vssd1
+ vccd1 vccd1 _00313_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11955_ _05799_ _05807_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__or2_2
XFILLER_0_118_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ _05157_ _05159_ _05161_ _05162_ _05163_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__a32o_2
XANTENNA__10210__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07685__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11886_ total_design.core.math.pc_val\[1\] total_design.core.program_count.imm_val_reg\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13625_ clknet_leaf_55_clk net1332 net1113 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10837_ _05090_ _05093_ _05095_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13556_ clknet_leaf_144_clk _01023_ net1181 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07437__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768_ _05026_ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09300__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12507_ net974 total_design.core.instr_mem.instruction_i\[17\] vssd1 vssd1 vccd1
+ vccd1 _01708_ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13487_ clknet_leaf_147_clk _00954_ net1152 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10699_ net265 net2808 net357 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12438_ net2765 net265 net347 vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12369_ _01622_ _01626_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14108_ clknet_leaf_99_clk _01288_ net1230 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07070__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14039_ clknet_leaf_83_clk _01219_ net1243 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[121\]
+ sky130_fd_sc_hd__dfrtp_1
X_06930_ total_design.core.regFile.register\[22\]\[7\] net776 net770 total_design.core.regFile.register\[7\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__a22o_1
XANTENNA__09898__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06861_ total_design.core.regFile.register\[0\]\[6\] net685 _02411_ _02417_ vssd1
+ vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_98_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08600_ total_design.data_in_BUS\[21\] net340 net714 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[21\]
+ sky130_fd_sc_hd__and3_1
X_09580_ _04105_ _04809_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__nand2_1
X_06792_ total_design.core.regFile.register\[21\]\[5\] net599 net568 total_design.core.regFile.register\[12\]\[5\]
+ _02350_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__a221o_1
X_14513__1285 vssd1 vssd1 vccd1 vccd1 net1285 _14513__1285/LO sky130_fd_sc_hd__conb_1
XFILLER_0_54_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08531_ _03879_ _03880_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08462_ _03787_ _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_102_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07413_ _02938_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__inv_2
X_08393_ net720 _03749_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[3\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_86_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07344_ total_design.core.regFile.register\[19\]\[15\] net825 _02872_ _02873_ vssd1
+ vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_154_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07428__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06393__X _01969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09210__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07275_ total_design.core.regFile.register\[2\]\[14\] net639 net570 total_design.core.regFile.register\[17\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06226_ _01798_ _01802_ _01804_ _01800_ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__and4bb_1
X_09014_ _04262_ _04266_ net467 vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06157_ total_design.core.regFile.register\[20\]\[0\] vssd1 vssd1 vccd1 vccd1 _01740_
+ sky130_fd_sc_hd__inv_2
Xhold120 total_design.core.data_mem.data_bus_i_reg\[19\] vssd1 vssd1 vccd1 vccd1 net1436
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 total_design.core.math.pc_val\[28\] vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1222_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold142 total_design.core.data_mem.data_read_adr_reg2\[18\] vssd1 vssd1 vccd1 vccd1
+ net1458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold153 total_design.core.data_mem.data_read_adr_reg2\[27\] vssd1 vssd1 vccd1 vccd1
+ net1469 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07061__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 total_design.core.data_mem.data_bus_i_reg\[23\] vssd1 vssd1 vccd1 vccd1 net1480
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 total_design.core.data_mem.data_cpu_i_reg\[26\] vssd1 vssd1 vccd1 vccd1 net1491
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07600__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold186 total_design.core.data_mem.data_read_adr_reg2\[14\] vssd1 vssd1 vccd1 vccd1
+ net1502 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A _02035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10803__B net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold197 total_design.lcd_display.row_1\[66\] vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 _02078_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_4
Xfanout611 _02072_ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__buf_4
Xfanout622 net623 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_8
X_09916_ _04118_ _04971_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__nor2_1
Xfanout633 _02061_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12488__A2 total_design.core.ctrl.instruction\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout644 _02056_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1108_X net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout655 net658 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__buf_6
Xfanout666 net669 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11696__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ net163 net2545 net437 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__mux2_1
Xfanout677 _02040_ vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__buf_4
Xfanout688 net689 vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_4
Xfanout699 net700 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ net168 net1898 net445 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__mux2_1
X_08729_ _00033_ _00031_ _00030_ _03987_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__nor4_1
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08313__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06728__B _02292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11740_ net1850 net956 _05049_ _05695_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10030__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08864__A1 total_design.core.ctrl.instruction\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_96_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06875__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout902_X net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11671_ _05613_ net1758 net129 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10818__X _05077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13410_ clknet_leaf_127_clk _00877_ net1192 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10622_ net171 net2481 net365 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__mux2_1
XANTENNA__08077__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14390_ clknet_leaf_197_clk _01531_ net1007 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11620__A0 _05477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13341_ clknet_leaf_14_clk _00808_ net1025 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10553_ net181 net1966 net375 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__mux2_1
XANTENNA__08092__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13960__RESET_B net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13272_ clknet_leaf_135_clk _00739_ net1187 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10484_ net193 net2566 net377 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__mux2_1
X_14537__1309 vssd1 vssd1 vccd1 vccd1 net1309 _14537__1309/LO sky130_fd_sc_hd__conb_1
X_12223_ total_design.core.math.pc_val\[9\] total_design.core.program_count.imm_val_reg\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07846__Y _03350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07052__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12154_ _06001_ _06004_ _06006_ _06008_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__or4_1
XANTENNA__11368__Y _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09592__A2 _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11105_ total_design.core.data_bus_o\[11\] _01728_ net515 net698 vssd1 vssd1 vccd1
+ vccd1 _05364_ sky130_fd_sc_hd__and4_1
XANTENNA__10205__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12085_ total_design.lcd_display.row_2\[68\] net349 _05832_ total_design.lcd_display.row_2\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11036_ net351 _05281_ _05285_ _05293_ _05279_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_21_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11384__X _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ clknet_leaf_149_clk _00454_ net1148 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11938_ _05798_ _05799_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__or2_2
XANTENNA__07658__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11869_ total_design.lcd_display.currentState\[3\] _05747_ total_design.lcd_display.currentState\[5\]
+ total_design.lcd_display.currentState\[4\] vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_60_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13608_ clknet_leaf_58_clk net1337 net1117 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08572__C net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09030__A _02182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11611__A0 _05648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13539_ clknet_leaf_16_clk _01006_ net1024 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08083__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07060_ total_design.core.regFile.register\[29\]\[10\] net655 net640 total_design.core.regFile.register\[19\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07830__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09684__B _04909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09583__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07962_ net553 total_design.core.data_mem.data_cpu_i\[27\] total_design.core.ctrl.imm_32\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10115__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08868__X _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11678__A0 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ _04925_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__inv_2
XANTENNA__09904__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06913_ _02453_ _02464_ _02465_ _02466_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_147_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07893_ total_design.core.regFile.register\[0\]\[26\] net875 _03394_ vssd1 vssd1
+ vccd1 vccd1 _03395_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ _04848_ _04859_ net450 vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_74_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06844_ total_design.core.regFile.register\[30\]\[6\] net661 net603 total_design.core.regFile.register\[31\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07897__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06829__A _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09205__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11454__B _05675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ _04710_ _04793_ net329 vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__mux2_1
X_06775_ net551 total_design.core.data_mem.data_cpu_i\[4\] _02336_ vssd1 vssd1 vccd1
+ vccd1 _02337_ sky130_fd_sc_hd__o21ai_4
XANTENNA__13723__Q total_design.core.data_cpu_o\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout263_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06548__B net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08514_ _03844_ _03850_ _03864_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_19_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_162_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09494_ _03134_ net447 _04366_ _04664_ _04727_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_121_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07649__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06857__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08445_ total_design.keypad0.key_out\[7\] _03753_ _03798_ vssd1 vssd1 vccd1 vccd1
+ _03799_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout430_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1172_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout149_X net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08763__B _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08376_ _01888_ _03733_ _03724_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__a21oi_1
Xwire308 _03015_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_4
XFILLER_0_163_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11602__A0 _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_177_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07327_ total_design.core.regFile.register\[28\]\[15\] net587 _02851_ _02856_ net688
+ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08074__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1058_X net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07282__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07258_ _02792_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout897_A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06209_ _01771_ _01787_ _01786_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_14_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09594__B _03322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07189_ total_design.core.regFile.register\[21\]\[12\] net761 _02727_ vssd1 vssd1
+ vccd1 vccd1 _02728_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10025__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout430 net433 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_6
Xfanout441 _04970_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11669__A0 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout452 _04121_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__buf_12
XPHY_EDGE_ROW_92_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout463 net464 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout852_X net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout474 _05805_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_6
Xfanout485 _05007_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__clkbuf_4
X_12910_ clknet_leaf_191_clk _00377_ net1032 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout496 net497 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_8
X_13890_ clknet_leaf_87_clk _01070_ net1250 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07888__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ clknet_leaf_177_clk _00308_ net1047 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12094__B1 _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12772_ clknet_leaf_106_clk _00239_ net1223 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14511_ net1283 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
X_11723_ _01731_ _01912_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__nand2_2
XANTENNA__06848__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10695__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11380__A _05612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14442_ clknet_leaf_61_clk net1358 net1216 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11654_ _05621_ net1678 net129 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10605_ net239 net2270 net366 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__mux2_1
X_14373_ clknet_leaf_171_clk _01514_ net1162 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11585_ _05630_ net1710 net144 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13324_ clknet_leaf_168_clk _00791_ net1156 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07273__B1 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10536_ net252 net2005 net376 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07812__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14512__1284 vssd1 vssd1 vccd1 vccd1 net1284 _14512__1284/LO sky130_fd_sc_hd__conb_1
XFILLER_0_122_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13255_ clknet_leaf_176_clk _00722_ net1048 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10467_ net274 net2066 net379 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__mux2_1
XANTENNA__10724__A total_design.core.instr_fetch vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12206_ _06037_ _06045_ _06046_ _06043_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_0_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07025__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13186_ clknet_leaf_131_clk _00653_ net1197 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10398_ net270 net2500 net387 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12137_ total_design.lcd_display.row_1\[95\] _05812_ _05838_ total_design.lcd_display.row_1\[31\]
+ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__a22o_1
XANTENNA__09009__B net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12068_ total_design.lcd_display.row_1\[115\] _05814_ _05829_ total_design.lcd_display.row_1\[107\]
+ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__a22o_1
XANTENNA__08848__B net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14247__RESET_B net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ _05275_ _05277_ _05055_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__a21o_2
XANTENNA__07879__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12085__B1 _05832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08289__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06560_ _01739_ total_design.core.regFile.register\[12\]\[1\] net918 _01948_ vssd1
+ vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__and4_1
XFILLER_0_87_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06839__B1 total_design.core.ctrl.instruction\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_47_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06491_ total_design.core.regFile.register\[14\]\[0\] net743 net730 net727 vssd1
+ vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__and4_1
XFILLER_0_129_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08230_ net1405 net544 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[13\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09031__Y _04283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08161_ net892 _02342_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[4\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08056__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07112_ total_design.core.regFile.register\[22\]\[11\] net677 net662 total_design.core.regFile.register\[30\]\[11\]
+ _02651_ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__a221o_1
X_08092_ total_design.core.regFile.register\[21\]\[30\] net599 net587 total_design.core.regFile.register\[28\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07803__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07043_ net751 _02589_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[9\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload40 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__inv_6
XFILLER_0_152_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload51 clknet_leaf_176_clk vssd1 vssd1 vccd1 vccd1 clkload51/X sky130_fd_sc_hd__clkbuf_8
Xclkload62 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_77_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload73 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 clkload73/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_77_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload84 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 clkload84/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__07016__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload95 clknet_leaf_147_clk vssd1 vssd1 vccd1 vccd1 clkload95/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13718__Q total_design.core.data_cpu_o\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07567__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08764__B1 _03350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08994_ net472 _03273_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1018_A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07945_ total_design.core.regFile.register\[8\]\[27\] net594 net563 total_design.core.regFile.register\[3\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__a22o_1
XANTENNA__06790__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08758__B _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07876_ total_design.core.regFile.register\[31\]\[26\] net832 net780 total_design.core.regFile.register\[27\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_3_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09615_ net186 net2551 net455 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__mux2_1
X_06827_ _02375_ _02377_ _02379_ _02386_ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__or4_2
XFILLER_0_74_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout645_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14536__1308 vssd1 vssd1 vccd1 vccd1 net1308 _14536__1308/LO sky130_fd_sc_hd__conb_1
XANTENNA__12076__B1 _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ total_design.core.math.pc_val\[21\] _04735_ total_design.core.math.pc_val\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__a21oi_1
X_06758_ total_design.core.regFile.register\[26\]\[4\] net644 net612 total_design.core.regFile.register\[11\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08295__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ net289 _04711_ _04707_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout812_A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__A1 _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06689_ total_design.core.regFile.register\[18\]\[3\] net860 net823 total_design.core.regFile.register\[19\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08428_ _03779_ _03780_ _03781_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload1 clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_136_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08359_ total_design.keypad0.key_out\[6\] total_design.keypad0.key_out\[7\] _03715_
+ _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__a211oi_1
XANTENNA__08047__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09809__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11370_ total_design.core.data_bus_o\[15\] net699 net510 vssd1 vssd1 vccd1 vccd1
+ _05629_ sky130_fd_sc_hd__a21o_1
X_10321_ net186 net1914 net493 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__mux2_1
XANTENNA__12473__A_N net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07007__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13040_ clknet_leaf_182_clk _00507_ net1040 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06233__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10252_ net198 net2216 net501 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__mux2_1
XANTENNA__06460__C net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ net172 net2358 net396 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__mux2_1
Xfanout1203 net1211 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__clkbuf_4
Xfanout1214 net1215 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08949__A total_design.core.ctrl.instruction\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1225 net1232 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__clkbuf_4
Xfanout1236 net1237 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__clkbuf_4
Xfanout1247 net1252 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input39_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1258 net1261 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout260 _04402_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_2
Xfanout271 _04348_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11375__A _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 net283 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_2
X_13942_ clknet_leaf_73_clk _01122_ net1209 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[88\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout293 _05696_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14459__Q total_design.core.instr_mem.instruction_adr_i\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13873_ clknet_leaf_68_clk total_design.core.ctrl.imm_32\[12\] net1111 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12824_ clknet_leaf_124_clk _00291_ net1186 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12755_ clknet_leaf_178_clk _00222_ net1035 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11706_ net10 net936 net879 net1847 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__a22o_1
X_12686_ clknet_leaf_189_clk _00153_ net1029 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14425_ clknet_leaf_29_clk total_design.core.data_out_INSTR\[20\] net1073 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11637_ _05657_ net1645 net135 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__mux2_1
XANTENNA__08038__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14356_ clknet_leaf_45_clk _00025_ net1086 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11568_ _05655_ net1711 net142 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13307_ clknet_leaf_143_clk _00774_ net1173 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold708 total_design.core.regFile.register\[15\]\[27\] vssd1 vssd1 vccd1 vccd1 net2024
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10519_ net186 net2096 net482 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__mux2_1
Xhold719 total_design.core.regFile.register\[4\]\[5\] vssd1 vssd1 vccd1 vccd1 net2035
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14287_ clknet_leaf_103_clk _01463_ net1238 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
X_11499_ net1531 _05670_ net151 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_139_Left_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13238_ clknet_leaf_155_clk _00705_ net1137 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06370__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08746__B1 _03206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13169_ clknet_leaf_148_clk _00636_ net1148 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08859__A total_design.core.ctrl.instruction\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1408 total_design.core.regFile.register\[2\]\[25\] vssd1 vssd1 vccd1 vccd1 net2724
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_144_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1419 total_design.core.regFile.register\[29\]\[23\] vssd1 vssd1 vccd1 vccd1 net2735
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06772__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ total_design.core.regFile.register\[3\]\[23\] net865 net842 total_design.core.regFile.register\[25\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__a22o_1
XANTENNA__09026__Y _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_140_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07661_ total_design.core.regFile.register\[26\]\[21\] net646 net590 total_design.core.regFile.register\[1\]\[21\]
+ _03171_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_140_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06524__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_148_Left_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09400_ _04617_ _04637_ _02941_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__a21oi_2
X_06612_ _02182_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__inv_2
XANTENNA__12058__B1 _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07592_ total_design.core.regFile.register\[10\]\[20\] net616 net608 total_design.core.regFile.register\[18\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09331_ _04221_ _04226_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__nand2_1
X_06543_ _02106_ net334 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07485__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09262_ _04416_ _04505_ net327 vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06474_ _01924_ net901 _02018_ total_design.core.ctrl.instruction\[18\] _01743_ vssd1
+ vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__o311a_1
XFILLER_0_28_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08213_ _03661_ _03663_ _03669_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_138_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08029__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09193_ _04439_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout226_A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08144_ _03628_ _03630_ _03632_ _03634_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__or4_2
XANTENNA__07237__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_157_Left_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload140 clknet_leaf_133_clk vssd1 vssd1 vccd1 vccd1 clkload140/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_116_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08075_ total_design.core.regFile.register\[27\]\[30\] net781 net766 total_design.core.regFile.register\[6\]\[30\]
+ _03568_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload151 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 clkload151/Y sky130_fd_sc_hd__inv_6
XANTENNA_fanout1135_A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06561__B net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload162 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 clkload162/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_113_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload173 clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 clkload173/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_3_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload184 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 clkload184/Y sky130_fd_sc_hd__clkinv_2
X_07026_ total_design.core.regFile.register\[29\]\[9\] net800 net785 total_design.core.regFile.register\[2\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout595_A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10544__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold13 total_design.core.data_mem.data_read_adr_reg\[18\] vssd1 vssd1 vccd1 vccd1
+ net1329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 total_design.core.data_mem.data_read_adr_reg\[7\] vssd1 vssd1 vccd1 vccd1
+ net1340 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _04227_ _04229_ net463 vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__mux2_1
XANTENNA__10811__B _05049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 total_design.core.math.pc_val\[13\] vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 total_design.core.data_mem.data_cpu_i_reg\[23\] vssd1 vssd1 vccd1 vccd1 net1362
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06763__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold57 total_design.core.math.pc_val\[14\] vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ total_design.core.regFile.register\[16\]\[27\] net855 net792 total_design.core.regFile.register\[24\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__a22o_1
XANTENNA__10303__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold68 total_design.core.math.pc_val\[18\] vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 total_design.core.data_mem.data_bus_i_reg\[29\] vssd1 vssd1 vccd1 vccd1 net1395
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__X _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_166_Left_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07859_ _03355_ _03357_ _03359_ _03361_ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14511__1283 vssd1 vssd1 vccd1 vccd1 net1283 _14511__1283/LO sky130_fd_sc_hd__conb_1
X_10870_ _05110_ _05128_ _05115_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__o21a_1
XANTENNA__06576__X total_design.core.data_mem.data_cpu_i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09529_ _03178_ _03180_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13733__RESET_B net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout815_X net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ net1427 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07476__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12471_ net2718 _01687_ _01689_ _01690_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14210_ clknet_leaf_60_clk _01390_ net1132 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11422_ net1643 _05624_ net159 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__mux2_1
XANTENNA__07228__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14141_ clknet_leaf_88_clk _01321_ net1258 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11353_ net303 _05608_ _05611_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_85_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10304_ net262 net2836 net494 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__mux2_1
X_14072_ clknet_leaf_109_clk _01252_ net1226 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[90\]
+ sky130_fd_sc_hd__dfrtp_1
X_11284_ _05484_ _05487_ _05542_ _05540_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__o31a_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13023_ clknet_leaf_182_clk _00490_ net1043 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10235_ net259 net2175 net502 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__mux2_1
XANTENNA__10535__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1011 net1014 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11376__Y _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07400__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1022 net1024 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_4
Xfanout1033 net1036 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__buf_2
X_10166_ net240 net2318 net397 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__mux2_1
XANTENNA__06754__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1044 net1045 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__buf_2
Xfanout1055 net1057 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_4
Xfanout1066 net1069 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__clkbuf_4
Xfanout1077 net1080 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__buf_2
XANTENNA__10213__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1088 net1089 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__clkbuf_4
X_10097_ net253 net2685 net402 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__mux2_1
Xfanout1099 net1104 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__buf_2
XFILLER_0_89_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13925_ clknet_leaf_85_clk _01105_ net1249 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11392__X _05651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload4_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13856_ clknet_leaf_56_clk _01064_ net1115 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08858__A_N total_design.core.ctrl.instruction\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12807_ clknet_leaf_176_clk _00274_ net1052 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08845__C _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13787_ clknet_leaf_57_clk total_design.core.data_mem.stored_data_adr\[30\] net1118
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[30\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10999_ _05250_ _05255_ _05244_ _05245_ _05247_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12738_ clknet_leaf_129_clk _00205_ net1198 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12669_ clknet_leaf_11_clk _00136_ net1020 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14408_ clknet_leaf_41_clk total_design.core.data_out_INSTR\[3\] net1090 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07219__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06190_ net998 net997 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_96_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_160_Right_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14339_ clknet_leaf_54_clk _01500_ net1110 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold505 net77 vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold516 total_design.data_in_BUS\[26\] vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 net99 vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 total_design.lcd_display.row_1\[97\] vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14535__1307 vssd1 vssd1 vccd1 vccd1 net1307 _14535__1307/LO sky130_fd_sc_hd__conb_1
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold549 total_design.core.math.pc_val\[2\] vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08900_ _02117_ _04153_ net459 vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__or3b_1
X_09880_ net166 net2387 net432 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _04079_ _04085_ _04033_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1205 total_design.core.regFile.register\[28\]\[6\] vssd1 vssd1 vccd1 vccd1 net2521
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 total_design.core.regFile.register\[11\]\[24\] vssd1 vssd1 vccd1 vccd1 net2532
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06745__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12279__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10123__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1227 total_design.core.regFile.register\[24\]\[2\] vssd1 vssd1 vccd1 vccd1 net2543
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ net307 _03322_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__nand2_1
Xhold1238 total_design.core.regFile.register\[31\]\[24\] vssd1 vssd1 vccd1 vccd1 net2554
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 total_design.core.regFile.register\[10\]\[12\] vssd1 vssd1 vccd1 vccd1 net2565
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07713_ _03215_ _03217_ _03219_ _03221_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__or4_1
XANTENNA__09912__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08693_ net1818 _03956_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout176_A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07644_ _03149_ _03155_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06837__A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07170__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13731__Q total_design.core.data_bus_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07575_ _01748_ _03041_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout343_A _01905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1085_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09314_ _02741_ net504 vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__or2_1
XANTENNA__07458__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06526_ total_design.core.regFile.register\[25\]\[0\] net647 _02069_ _02071_ _02077_
+ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_91_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09245_ _02587_ net504 net446 _02585_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout131_X net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06457_ _01923_ net896 _02019_ _01745_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1252_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07668__A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09176_ total_design.core.math.pc_val\[6\] _04397_ vssd1 vssd1 vccd1 vccd1 _04424_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06388_ net926 net948 net912 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08127_ total_design.core.regFile.register\[18\]\[31\] net858 net781 total_design.core.regFile.register\[27\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07630__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08058_ net306 _03552_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06984__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10780__A3 total_design.core.data_bus_o\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07009_ total_design.core.regFile.register\[1\]\[9\] net590 net575 total_design.core.regFile.register\[24\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__a22o_1
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__clkbuf_4
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__clkbuf_4
X_10020_ net286 net1969 net413 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06736__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10033__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__A2_N net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08011__B _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09822__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ _05746_ _05749_ _05807_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__or3_2
XANTENNA__08489__A2 _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13710_ clknet_leaf_32_clk total_design.core.data_mem.stored_read_data\[17\] net1063
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[17\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11493__A1 _05626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10922_ _05157_ _05159_ _05155_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__a21o_1
XANTENNA__07161__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13641_ clknet_leaf_55_clk total_design.core.data_mem.data_write_adr_i\[13\] net1117
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[13\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11372__B _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10853_ _05095_ _05099_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07449__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13572_ clknet_leaf_38_clk total_design.core.data_mem.data_bus_i\[8\] net1078 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[8\] sky130_fd_sc_hd__dfrtp_1
X_10784_ total_design.core.data_bus_o\[18\] net696 _05042_ net517 vssd1 vssd1 vccd1
+ vccd1 _05043_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_82_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12523_ net975 total_design.core.instr_mem.instruction_i\[25\] vssd1 vssd1 vccd1
+ vccd1 _01716_ sky130_fd_sc_hd__and2b_1
XFILLER_0_87_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12454_ net1960 net195 net344 vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11405_ _05077_ _05610_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__nor2_1
X_12385_ net991 _01643_ _01644_ _01645_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_10_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10208__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14124_ clknet_leaf_99_clk _01304_ net1230 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11336_ _05529_ _05536_ _05534_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11387__X _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06975__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14055_ clknet_leaf_83_clk _01235_ net1241 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[73\]
+ sky130_fd_sc_hd__dfrtp_1
X_11267_ _05514_ _05517_ _05518_ _05519_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_24_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13006_ clknet_leaf_187_clk _00473_ net1031 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10218_ _04842_ net2540 net391 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__mux2_1
X_11198_ total_design.core.data_bus_o\[18\] net695 net510 vssd1 vssd1 vccd1 vccd1
+ _05457_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10149_ net173 net2796 net401 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11484__A1 _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13908_ clknet_leaf_111_clk _01088_ net1209 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07688__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08575__C net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13839_ clknet_leaf_59_clk _01047_ net1126 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07360_ net552 total_design.core.data_mem.data_cpu_i\[15\] total_design.core.ctrl.imm_32\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06944__X total_design.core.ctrl.imm_32\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06311_ _01808_ _01840_ _01841_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_21_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07291_ total_design.core.regFile.register\[24\]\[14\] net793 _02822_ _02823_ vssd1
+ vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_135_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11502__S net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09179__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09030_ _02182_ net462 vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__and2_1
X_06242_ net961 _01820_ _01819_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07860__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06173_ total_design.core.data_cpu_o\[8\] vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__inv_2
XANTENNA__10118__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold302 total_design.lcd_display.row_2\[54\] vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold313 total_design.lcd_display.row_2\[77\] vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 total_design.lcd_display.row_1\[29\] vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07612__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09907__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold335 total_design.lcd_display.row_2\[50\] vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 total_design.lcd_display.row_2\[101\] vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 total_design.lcd_display.row_2\[37\] vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold368 total_design.lcd_display.row_1\[90\] vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ net235 net2806 net425 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__mux2_1
Xhold379 total_design.lcd_display.row_1\[122\] vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout804 net805 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout815 _01969_ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09365__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout826 _01964_ vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__buf_4
X_09863_ net228 net2745 net430 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__mux2_1
Xfanout837 _01958_ vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_4
Xfanout848 net849 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_4
XANTENNA__06718__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net860 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__buf_4
Xhold1002 total_design.core.regFile.register\[17\]\[11\] vssd1 vssd1 vccd1 vccd1 net2318
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08814_ total_design.core.data_mem.data_cpu_i\[2\] _02233_ vssd1 vssd1 vccd1 vccd1
+ _04069_ sky130_fd_sc_hd__or2_1
Xhold1013 total_design.core.regFile.register\[27\]\[4\] vssd1 vssd1 vccd1 vccd1 net2329
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 total_design.core.regFile.register\[30\]\[26\] vssd1 vssd1 vccd1 vccd1 net2340
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ net230 net2245 net438 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__mux2_1
Xhold1035 total_design.core.regFile.register\[2\]\[19\] vssd1 vssd1 vccd1 vccd1 net2351
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 total_design.core.regFile.register\[30\]\[28\] vssd1 vssd1 vccd1 vccd1 net2362
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1057 total_design.core.regFile.register\[6\]\[16\] vssd1 vssd1 vccd1 vccd1 net2373
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ _03064_ _03083_ _03112_ net457 vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__o22a_1
Xhold1068 total_design.core.regFile.register\[4\]\[31\] vssd1 vssd1 vccd1 vccd1 net2384
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 total_design.core.regFile.register\[19\]\[12\] vssd1 vssd1 vccd1 vccd1 net2395
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12121__C1 _05971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_X net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__A1 _05636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07679__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08676_ total_design.keypad0.counter\[6\] total_design.keypad0.counter\[7\] _03952_
+ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_159_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11192__B _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07627_ total_design.core.regFile.register\[10\]\[21\] net836 net791 total_design.core.regFile.register\[24\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07558_ total_design.core.regFile.register\[26\]\[19\] net870 net784 total_design.core.regFile.register\[2\]\[19\]
+ _03075_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08782__A _02565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06509_ net744 net738 net726 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07489_ total_design.core.regFile.register\[7\]\[18\] net651 _03009_ net686 vssd1
+ vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__a211o_1
XFILLER_0_174_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09228_ _01755_ net752 _04473_ net905 _04470_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__o221a_2
XANTENNA__06654__A1 total_design.core.regFile.register\[29\]\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07851__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09159_ _02442_ net703 _04406_ net533 vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__a211o_1
XANTENNA__10028__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09817__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ _06012_ _06015_ _06020_ _06021_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__a211oi_1
XANTENNA__07603__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06957__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ net515 _05094_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__nand2_2
Xhold880 total_design.core.regFile.register\[19\]\[22\] vssd1 vssd1 vccd1 vccd1 net2196
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold891 total_design.core.regFile.register\[26\]\[3\] vssd1 vssd1 vccd1 vccd1 net2207
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06241__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11052_ _05306_ _05307_ _05308_ _05310_ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__or4_1
XANTENNA__06709__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ _04681_ net2162 net414 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__mux2_1
XANTENNA__11702__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09552__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07382__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11466__A1 _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09124__Y _04374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11954_ _05803_ _05807_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_28_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07134__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10905_ _05162_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_28_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14534__1306 vssd1 vssd1 vccd1 vccd1 net1306 _14534__1306/LO sky130_fd_sc_hd__conb_1
X_11885_ total_design.core.math.pc_val\[1\] total_design.core.program_count.imm_val_reg\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_192_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_192_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_103_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13624_ clknet_leaf_56_clk net1342 net1113 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10836_ net521 _05094_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__nand2_2
XFILLER_0_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13555_ clknet_leaf_180_clk _01022_ net1042 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08095__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10767_ _01859_ _01869_ _01887_ _05025_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_41_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12506_ net976 total_design.core.ctrl.instruction\[16\] net881 _01707_ vssd1 vssd1
+ vccd1 vccd1 _01555_ sky130_fd_sc_hd__a22o_1
XANTENNA__07842__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__B _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13486_ clknet_leaf_188_clk _00953_ net1029 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10698_ net273 net2529 net360 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12437_ net1936 net272 net346 vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09727__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12368_ _01630_ total_design.core.math.pc_val\[24\] net523 vssd1 vssd1 vccd1 vccd1
+ _01494_ sky130_fd_sc_hd__mux2_1
XANTENNA__06940__A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06948__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14107_ clknet_leaf_90_clk _01287_ net1260 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_112_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11319_ net294 _05568_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12299_ net992 _06134_ _06135_ _06136_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_39_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14038_ clknet_leaf_100_clk _01218_ net1229 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09028__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06860_ _02413_ _02414_ _02415_ _02416_ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__or4_1
XFILLER_0_101_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06939__X _02492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07373__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__A _03273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06791_ total_design.core.regFile.register\[30\]\[5\] net661 net610 total_design.core.regFile.register\[18\]\[5\]
+ _02349_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08530_ _03866_ _03878_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__nand2_1
XANTENNA__11457__A1 _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10401__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_121_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07125__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08461_ _03813_ _03814_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_183_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_183_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07412_ _02917_ _02937_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08392_ total_design.data_in_BUS\[3\] _01905_ _03748_ vssd1 vssd1 vccd1 vccd1 _03749_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_102_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08086__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07343_ total_design.core.regFile.register\[18\]\[15\] net858 net785 total_design.core.regFile.register\[2\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout139_A _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07833__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07274_ total_design.core.regFile.register\[21\]\[14\] net600 net596 total_design.core.regFile.register\[8\]\[14\]
+ _02806_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09013_ _04265_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_171_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06225_ total_design.core.data_adr_o\[28\] _01803_ net961 vssd1 vssd1 vccd1 vccd1
+ _01804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1048_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 total_design.core.instr_mem.instruction_adr_stored\[11\] vssd1 vssd1 vccd1
+ vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold121 total_design.core.instr_mem.instruction_adr_stored\[21\] vssd1 vssd1 vccd1
+ vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
X_06156_ total_design.core.ctrl.instruction\[24\] vssd1 vssd1 vccd1 vccd1 _01739_
+ sky130_fd_sc_hd__inv_2
Xhold132 total_design.core.instr_mem.instruction_adr_stored\[25\] vssd1 vssd1 vccd1
+ vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 total_design.core.instr_mem.instruction_adr_stored\[24\] vssd1 vssd1 vccd1
+ vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold154 total_design.core.data_mem.data_read_adr_reg2\[22\] vssd1 vssd1 vccd1 vccd1
+ net1470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold165 total_design.core.data_mem.data_read_adr_reg2\[12\] vssd1 vssd1 vccd1 vccd1
+ net1481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 total_design.core.data_mem.data_read_adr_reg2\[1\] vssd1 vssd1 vccd1 vccd1
+ net1492 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1215_A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold187 net53 vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _02076_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09338__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold198 total_design.lcd_display.row_2\[97\] vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 net615 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__clkbuf_8
X_09915_ net164 net2022 net428 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__mux2_1
Xfanout623 _02066_ vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_4
Xfanout634 _02061_ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout675_A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 net646 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout656 net658 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_8
Xfanout667 net669 vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_8
X_09846_ net167 net2665 net436 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__mux2_1
Xfanout678 net681 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__clkbuf_8
Xfanout689 _02034_ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09777_ net170 net2492 net442 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__mux2_1
X_06989_ _02536_ _02538_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_126_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout842_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08728_ _03971_ _00035_ _00036_ _03986_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__or4_1
XANTENNA__11448__A1 _05645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10311__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06297__A _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07116__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11999__A2 _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08659_ _03941_ net711 _03940_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__and3b_1
XFILLER_0_139_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_174_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_174_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08864__A2 total_design.core.ctrl.instruction\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11670_ _05657_ net1699 net130 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10621_ net172 net2290 net367 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__mux2_1
XANTENNA__08077__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13340_ clknet_leaf_12_clk _00807_ net1026 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10552_ net188 net2215 net375 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06236__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13271_ clknet_leaf_124_clk _00738_ net1186 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10483_ net199 net2138 net378 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12222_ _06062_ _06063_ _06060_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ total_design.lcd_display.row_2\[47\] _05844_ _05846_ total_design.lcd_display.row_2\[103\]
+ _06007_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11104_ total_design.core.data_bus_o\[11\] _05049_ _05059_ _05064_ net515 vssd1 vssd1
+ vccd1 vccd1 _05363_ sky130_fd_sc_hd__o2111a_1
XANTENNA__11097__B _05220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12084_ total_design.lcd_display.row_2\[44\] _05844_ _05845_ total_design.lcd_display.row_2\[20\]
+ _05941_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11035_ net351 _05281_ _05285_ _05293_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__a211oi_1
XANTENNA__08001__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07355__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12986_ clknet_leaf_124_clk _00453_ net1188 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07107__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12100__A2 _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14197__Q net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11937_ _05745_ _05749_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_165_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_165_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07512__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08855__A2 _04102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11868_ total_design.lcd_display.currentState\[4\] _05747_ vssd1 vssd1 vccd1 vccd1
+ _05751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09311__A _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13607_ clknet_leaf_62_clk net1345 net1125 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10819_ total_design.core.data_bus_o\[9\] net698 vssd1 vssd1 vccd1 vccd1 _05078_
+ sky130_fd_sc_hd__nand2_2
XANTENNA__08068__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11799_ total_design.lcd_display.cnt_20ms\[0\] total_design.lcd_display.cnt_20ms\[1\]
+ net2163 vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07815__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13538_ clknet_leaf_126_clk _01005_ net1193 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13469_ clknet_leaf_9_clk _00936_ net1020 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08214__X total_design.core.data_mem.next_write vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06670__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07961_ net553 total_design.core.data_mem.data_cpu_i\[27\] total_design.core.ctrl.imm_32\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__a21o_1
XANTENNA__13670__RESET_B net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ total_design.core.math.pc_val\[29\] _04905_ vssd1 vssd1 vccd1 vccd1 _04925_
+ sky130_fd_sc_hd__xnor2_1
X_06912_ total_design.core.regFile.register\[20\]\[7\] net673 net569 total_design.core.regFile.register\[17\]\[7\]
+ _02451_ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__a221o_1
X_07892_ total_design.core.regFile.register\[17\]\[26\] net820 _03377_ _03380_ _03393_
+ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_147_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07346__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ net314 net296 _04296_ _04849_ _04858_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__o311a_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09740__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06843_ total_design.core.regFile.register\[2\]\[6\] net638 net622 total_design.core.regFile.register\[4\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10131__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09562_ net468 _04749_ _04792_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11454__C _05478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09205__B _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06774_ net555 total_design.core.ctrl.imm_32\[4\] vssd1 vssd1 vccd1 vccd1 _02336_
+ sky130_fd_sc_hd__or2_1
X_08513_ _03861_ _03863_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__nor2_1
XANTENNA__09920__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09493_ net968 _03134_ _03135_ net537 vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_78_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09699__Y _04924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_156_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_156_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout256_A _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08444_ _03797_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08375_ total_design.keypad0.key_out\[2\] _03732_ _03719_ vssd1 vssd1 vccd1 vccd1
+ _03733_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout423_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire309 _02988_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_4
XFILLER_0_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07326_ total_design.core.regFile.register\[29\]\[15\] net657 net645 total_design.core.regFile.register\[26\]\[15\]
+ _02855_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07257_ _02770_ _02789_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_30_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12158__A2 _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06208_ total_design.core.instr_mem.instruction_adr_i\[9\] total_design.core.instr_mem.instruction_adr_stored\[9\]
+ net984 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07188_ total_design.core.regFile.register\[31\]\[12\] net833 net788 total_design.core.regFile.register\[13\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout792_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1120_X net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10306__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14533__1305 vssd1 vssd1 vccd1 vccd1 net1305 _14533__1305/LO sky130_fd_sc_hd__conb_1
XFILLER_0_2_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07585__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06793__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout420 net421 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_4
Xfanout431 net433 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_6
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout442 _04969_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_6
Xfanout453 _04117_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13340__RESET_B net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout464 _02184_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_2
Xfanout475 _05797_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_2
XANTENNA__07337__A2 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout486 _05007_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_6_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09829_ net230 net1905 net434 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__mux2_1
Xfanout497 _05004_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_4
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10041__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ clknet_leaf_24_clk _00307_ net1108 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09830__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12771_ clknet_leaf_6_clk _00238_ net1017 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_147_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_147_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11722_ net1507 net956 _05692_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__a21bo_1
X_14510_ net72 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_81_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11380__B _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14441_ clknet_leaf_64_clk net1865 net1134 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11653_ _05477_ net1831 net129 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11054__C1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10604_ net241 net2060 net368 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__mux2_1
X_14372_ clknet_leaf_177_clk _01513_ net1047 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11584_ _05651_ net1813 net141 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13323_ clknet_leaf_120_clk _00790_ net1191 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10535_ net264 net2761 net376 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11600__S net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12149__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09277__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13254_ clknet_leaf_200_clk _00721_ net1001 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10466_ net258 net2514 net379 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10724__B net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12205_ _06051_ _06052_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__nand2_1
XANTENNA__14480__Q total_design.core.ctrl.instruction\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_122_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10216__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13185_ clknet_leaf_123_clk _00652_ net1167 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10397_ net279 net2018 net387 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12136_ total_design.lcd_display.row_1\[47\] _05821_ _05841_ total_design.lcd_display.row_1\[15\]
+ _05990_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12067_ _05920_ _05922_ _05923_ _05925_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_53_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12431__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07328__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11018_ _05276_ _05255_ _05250_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__mux2_1
XANTENNA__13824__Q total_design.core.data_access vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06368__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08289__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_138_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_138_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12969_ clknet_leaf_17_clk _00436_ net1046 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06490_ net741 net730 net726 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07500__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08160_ net892 _02292_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07111_ total_design.core.regFile.register\[29\]\[11\] net658 _02092_ total_design.core.regFile.register\[12\]\[11\]
+ _02652_ vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07264__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08091_ total_design.core.regFile.register\[24\]\[30\] net575 _03581_ _03583_ net688
+ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_125_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11510__S net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload30 clknet_leaf_184_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__clkinv_4
X_07042_ _02544_ _02588_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__xor2_2
XFILLER_0_3_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload41 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__bufinv_16
Xclkload52 clknet_leaf_177_clk vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_77_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload63 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__clkinv_8
Xclkload74 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__inv_8
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload85 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload96 clknet_leaf_148_clk vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__inv_6
XANTENNA__10126__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10020__A0 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07567__A2 total_design.core.data_mem.data_cpu_i\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08764__A1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06550__D net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08764__B2 _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ net297 _04245_ _04217_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07944_ total_design.core.regFile.register\[20\]\[27\] net671 net571 total_design.core.regFile.register\[17\]\[27\]
+ _03442_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_166_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07875_ total_design.core.regFile.register\[29\]\[26\] net799 net760 total_design.core.regFile.register\[21\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_3_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout373_A _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09614_ net507 _04842_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__and2_1
X_06826_ total_design.core.regFile.register\[13\]\[5\] net788 _02381_ _02382_ _02385_
+ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_168_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09545_ total_design.core.math.pc_val\[21\] total_design.core.math.pc_val\[22\] _04735_
+ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06757_ total_design.core.regFile.register\[21\]\[4\] net597 net589 total_design.core.regFile.register\[1\]\[4\]
+ _02317_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_129_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout540_A _03676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_174_Right_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09476_ _04622_ _04709_ net329 vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__mux2_1
X_06688_ total_design.core.regFile.register\[12\]\[3\] net774 net772 total_design.core.regFile.register\[28\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__a22o_1
XANTENNA__06575__A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08427_ total_design.keypad0.key_out\[11\] total_design.keypad0.key_out\[8\] vssd1
+ vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout805_A _01974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08358_ net933 total_design.keypad0.key_out\[10\] total_design.keypad0.key_out\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload2 clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__inv_8
XANTENNA__11587__A0 _05477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07309_ _02839_ _02840_ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__or2_1
X_08289_ total_design.core.data_mem.data_write_adr_reg\[2\] net549 net540 total_design.core.data_mem.data_read_adr_reg\[2\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11420__S net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10320_ net189 net2625 net493 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06463__C1 total_design.core.ctrl.instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_131_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10251_ net201 net2680 net501 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__mux2_1
XANTENNA__10036__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07558__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09825__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08755__A1 _02968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ net176 net2282 net395 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__mux2_1
XANTENNA__06766__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1204 net1211 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__clkbuf_2
Xfanout1215 net1222 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__clkbuf_2
Xfanout1226 net1232 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__clkbuf_2
Xfanout1237 net1240 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__clkbuf_4
Xfanout250 net252 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1248 net1252 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__buf_2
Xfanout1259 net1261 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout261 net264 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout272 net275 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_2
X_13941_ clknet_leaf_92_clk _01121_ net1262 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[87\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout283 _04374_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_2
Xfanout294 _05463_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07715__C1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06469__B net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13872_ clknet_leaf_68_clk total_design.core.ctrl.imm_32\[11\] net1111 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07730__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12823_ clknet_leaf_163_clk _00290_ net1164 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12754_ clknet_leaf_137_clk _00221_ net1184 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11705_ net9 net934 net877 net2217 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__o22a_1
X_12685_ clknet_leaf_3_clk _00152_ net1011 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11636_ _05671_ net1700 net134 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__mux2_1
X_14424_ clknet_leaf_37_clk total_design.core.data_out_INSTR\[19\] net1076 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[19\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06772__X _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11578__A0 _05648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14355_ clknet_leaf_45_clk _00024_ net1086 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11567_ _05679_ net1760 net143 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10518_ net190 net2219 net482 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__mux2_1
X_13306_ clknet_leaf_134_clk _00773_ net1189 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14286_ net987 _01462_ net1082 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_12_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold709 total_design.core.regFile.register\[31\]\[4\] vssd1 vssd1 vccd1 vccd1 net2025
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11498_ net1598 _05667_ net149 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12860__CLK clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13237_ clknet_leaf_157_clk _00704_ net1141 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08787__A_N _02770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10449_ net203 net2328 net382 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07549__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_161_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08746__A1 _03157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06370__D net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08746__B2 _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13168_ clknet_leaf_186_clk _00635_ net1038 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06757__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08859__B total_design.core.ctrl.instruction\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11750__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ total_design.lcd_display.row_1\[54\] _05840_ _05848_ total_design.lcd_display.row_2\[126\]
+ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13099_ clknet_leaf_114_clk _00566_ net1202 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1409 total_design.core.regFile.register\[5\]\[29\] vssd1 vssd1 vccd1 vccd1 net2725
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_144_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_176_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07660_ total_design.core.regFile.register\[23\]\[21\] net679 net618 total_design.core.regFile.register\[10\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_140_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07182__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06611_ _02178_ _02180_ _02181_ _02152_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__o31a_4
X_07591_ total_design.core.regFile.register\[13\]\[20\] net666 net562 total_design.core.regFile.register\[3\]\[20\]
+ _03104_ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ _02796_ net701 _04570_ net533 vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__a211o_1
XFILLER_0_172_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06542_ _02106_ net470 vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__nand2b_4
X_14532__1304 vssd1 vssd1 vccd1 vccd1 net1304 _14532__1304/LO sky130_fd_sc_hd__conb_1
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09261_ _04458_ _04503_ net460 vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__mux2_1
X_06473_ total_design.core.regFile.register\[13\]\[0\] _02031_ net729 net727 vssd1
+ vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__and4_1
X_08212_ _03666_ _03668_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09192_ _04237_ _04241_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__or2_1
XANTENNA__11569__A0 _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08143_ total_design.core.regFile.register\[16\]\[31\] net634 net578 total_design.core.regFile.register\[27\]\[31\]
+ _03633_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout219_A _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07788__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload130 clknet_leaf_145_clk vssd1 vssd1 vccd1 vccd1 clkload130/Y sky130_fd_sc_hd__clkinv_2
X_08074_ total_design.core.regFile.register\[14\]\[30\] net863 net825 total_design.core.regFile.register\[19\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload141 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 clkload141/Y sky130_fd_sc_hd__clkinv_4
Xclkload152 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 clkload152/Y sky130_fd_sc_hd__inv_8
XANTENNA__06561__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload163 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 clkload163/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_168_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07025_ total_design.core.regFile.register\[31\]\[9\] net833 net769 total_design.core.regFile.register\[7\]\[9\]
+ _02572_ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a221o_1
Xclkload174 clknet_leaf_87_clk vssd1 vssd1 vccd1 vccd1 clkload174/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_168_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_129_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1128_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout490_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__B1 _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08769__B net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 total_design.core.data_mem.data_read_adr_reg\[13\] vssd1 vssd1 vccd1 vccd1
+ net1330 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ net473 _02564_ _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__o21ai_1
Xhold25 total_design.core.data_mem.data_read_adr_reg\[15\] vssd1 vssd1 vccd1 vccd1
+ net1341 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10811__C _05064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold36 total_design.core.data_mem.data_bus_i_reg\[0\] vssd1 vssd1 vccd1 vccd1 net1352
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 total_design.core.data_mem.data_cpu_i_reg\[11\] vssd1 vssd1 vccd1 vccd1 net1363
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold58 total_design.core.data_mem.data_cpu_i_reg\[22\] vssd1 vssd1 vccd1 vccd1 net1374
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ total_design.core.regFile.register\[30\]\[27\] net839 net811 total_design.core.regFile.register\[23\]\[27\]
+ _03423_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__a221o_1
Xhold69 total_design.core.data_mem.data_cpu_i_reg\[29\] vssd1 vssd1 vccd1 vccd1 net1385
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout755_A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09162__A1 _04409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ total_design.core.regFile.register\[11\]\[25\] net613 net609 total_design.core.regFile.register\[18\]\[25\]
+ _03360_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07173__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07712__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12049__A1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06809_ total_design.core.regFile.register\[25\]\[5\] net844 net833 total_design.core.regFile.register\[31\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07789_ total_design.core.regFile.register\[27\]\[24\] net780 net768 total_design.core.regFile.register\[7\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout922_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06920__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09528_ net203 net1987 net455 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09459_ _04685_ _04686_ _04694_ net449 vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout808_X net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12470_ total_design.keypad0.key_counter\[2\] _01687_ vssd1 vssd1 vccd1 vccd1 _01690_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11421_ net1593 _05635_ net158 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07779__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14140_ clknet_leaf_109_clk _01320_ net1228 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11352_ net514 _05035_ _05459_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10303_ net266 net2541 net492 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__mux2_1
X_14071_ clknet_leaf_84_clk _01251_ net1245 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11283_ _05498_ _05504_ _05541_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13022_ clknet_leaf_175_clk _00489_ net1053 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12524__A2 total_design.core.ctrl.instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10234_ net281 net1911 net500 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__mux2_1
Xfanout1001 net1002 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_4
Xfanout1012 net1014 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_4
X_10165_ net254 net2563 net394 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__mux2_1
Xfanout1023 net1024 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_4
Xfanout1034 net1036 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1045 net1059 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__buf_2
XANTENNA__07951__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1056 net1057 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__clkbuf_4
X_10096_ net249 net2520 net403 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__mux2_1
Xfanout1067 net1069 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__buf_2
Xfanout1078 net1080 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09689__C1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1089 net1105 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13924_ clknet_leaf_97_clk _01104_ net1244 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07164__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07703__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13855_ clknet_leaf_57_clk _01063_ net1118 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06911__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ clknet_leaf_201_clk _00273_ net1003 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13786_ clknet_leaf_55_clk total_design.core.data_mem.stored_data_adr\[29\] net1117
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[29\] sky130_fd_sc_hd__dfrtp_1
X_10998_ _05227_ _05244_ _05234_ _05228_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_48_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07104__A _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12737_ clknet_leaf_122_clk _00204_ net1169 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07598__X _03112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12668_ clknet_leaf_29_clk _00135_ net1073 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14407_ clknet_leaf_40_clk total_design.core.data_out_INSTR\[2\] net1092 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11619_ _05478_ _05480_ _05674_ _05675_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__or4_4
XFILLER_0_143_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06690__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10223__A0 _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12599_ clknet_leaf_161_clk _00066_ net1164 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14338_ clknet_leaf_53_clk _01499_ net1109 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[29\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold506 total_design.lcd_display.row_2\[4\] vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06978__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold517 total_design.lcd_display.row_1\[1\] vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06381__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold528 total_design.lcd_display.cnt_20ms\[10\] vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 total_design.core.regFile.register\[27\]\[1\] vssd1 vssd1 vccd1 vccd1 net1855
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14269_ clknet_leaf_47_clk _00001_ net1098 vssd1 vssd1 vccd1 vccd1 wishbone.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_111_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09392__A1 _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08830_ _04035_ _04044_ _04084_ _04045_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__a31o_1
XANTENNA__10404__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1206 total_design.keypad0.counter\[15\] vssd1 vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07942__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1217 total_design.core.regFile.register\[1\]\[2\] vssd1 vssd1 vccd1 vccd1 net2533
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08761_ _03395_ _03415_ _03440_ _03459_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__o22a_1
Xhold1228 total_design.core.regFile.register\[27\]\[18\] vssd1 vssd1 vccd1 vccd1 net2544
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 total_design.core.regFile.register\[25\]\[16\] vssd1 vssd1 vccd1 vccd1 net2555
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09144__A1 _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07712_ total_design.core.regFile.register\[11\]\[22\] net613 net574 total_design.core.regFile.register\[24\]\[22\]
+ _03220_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08692_ _03957_ _03964_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__nor2_1
X_07643_ total_design.core.regFile.register\[2\]\[21\] net784 _03151_ _03152_ _03154_
+ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06902__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06837__B _02395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07574_ net749 _03090_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[19\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06556__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09313_ net316 _04361_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__nand2_1
X_06525_ total_design.core.regFile.register\[8\]\[0\] net593 _02084_ _02051_ _02059_
+ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout336_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_146_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09244_ net313 _04275_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_157_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06456_ _01924_ net901 _02018_ total_design.core.ctrl.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 _02030_ sky130_fd_sc_hd__o31a_1
XFILLER_0_173_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09175_ _04407_ _04414_ _04422_ net450 vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__a31o_1
XANTENNA__07668__B total_design.core.ctrl.imm_32\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06681__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06387_ _01738_ net965 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout503_A _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ total_design.core.regFile.register\[25\]\[31\] net843 _03616_ _03617_ vssd1
+ vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__a211o_1
XFILLER_0_160_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06433__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08057_ net553 total_design.core.data_mem.data_cpu_i\[29\] total_design.core.ctrl.imm_32\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07008_ total_design.core.regFile.register\[9\]\[9\] net665 net657 total_design.core.regFile.register\[29\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__a22o_1
XANTENNA__09228__X _04474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10780__A4 total_design.core.data_bus_o\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10314__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1200_X net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07394__B1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ _02114_ _04211_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11970_ net531 _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__nor2_4
XANTENNA__07146__B1 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10921_ _05164_ _05179_ _05165_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__a21boi_2
XANTENNA_fanout925_X net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13640_ clknet_leaf_58_clk total_design.core.data_mem.data_write_adr_i\[12\] net1117
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[12\] sky130_fd_sc_hd__dfrtp_1
X_10852_ net521 _05048_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__nand2_2
XFILLER_0_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06466__C net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10783_ _05038_ _05039_ _05040_ _05041_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__or4_2
X_13571_ clknet_leaf_42_clk total_design.core.data_mem.data_bus_i\[7\] net1084 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[7\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_51_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12522_ net974 total_design.core.ctrl.instruction\[24\] net881 _01715_ vssd1 vssd1
+ vccd1 vccd1 _01563_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12453_ total_design.core.regFile.register\[31\]\[22\] net197 net345 vssd1 vssd1
+ vccd1 vccd1 _01524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10205__A0 _04588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06482__B net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ net302 _05653_ _05661_ _05662_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_151_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12384_ net991 _04863_ net894 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14123_ clknet_leaf_88_clk _01303_ net1251 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11335_ _05591_ _05592_ _05463_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_91_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11266_ _05516_ _05522_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__xnor2_1
X_14054_ clknet_leaf_100_clk _01234_ net1236 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10732__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09374__A1 total_design.core.data_cpu_o\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10217_ net189 net2479 net391 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__mux2_1
X_13005_ clknet_leaf_0_clk _00472_ net1003 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14531__1303 vssd1 vssd1 vccd1 vccd1 net1303 _14531__1303/LO sky130_fd_sc_hd__conb_1
XANTENNA__10224__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11197_ _05450_ _05455_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07924__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ net178 net2169 net401 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10079_ net187 net2469 net407 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07137__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12130__B1 _05814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ clknet_leaf_90_clk _01087_ net1263 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13838_ clknet_leaf_54_clk _01046_ net1109 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13769_ clknet_leaf_58_clk total_design.core.data_mem.stored_data_adr\[12\] net1126
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[12\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_42_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06310_ _01808_ _01843_ _01844_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__or3_1
XANTENNA__08101__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07290_ total_design.core.regFile.register\[9\]\[14\] net850 net818 total_design.core.regFile.register\[20\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__a22o_1
XANTENNA__06673__A _02213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06241_ total_design.core.instr_mem.instruction_adr_i\[31\] total_design.core.instr_mem.instruction_adr_stored\[31\]
+ net983 vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06172_ total_design.core.data_cpu_o\[7\] vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09062__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold303 total_design.lcd_display.row_1\[53\] vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold314 total_design.lcd_display.row_1\[101\] vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07775__Y _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold325 total_design.lcd_display.row_2\[74\] vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold336 total_design.lcd_display.row_2\[52\] vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold347 total_design.lcd_display.row_2\[103\] vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold358 total_design.lcd_display.row_2\[102\] vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 total_design.lcd_display.row_2\[69\] vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ net228 net2695 net422 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_3__f_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__06820__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout805 _01974_ vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_4
XFILLER_0_68_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout816 net818 vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_4_7__f_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14412__RESET_B net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10134__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09862_ net239 net2094 net432 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__mux2_1
Xfanout827 net830 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_8
Xfanout838 net841 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_8
Xfanout849 _01953_ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__buf_4
XANTENNA__07376__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09923__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1003 total_design.core.regFile.register\[27\]\[21\] vssd1 vssd1 vccd1 vccd1 net2319
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ _04067_ _04065_ _04064_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__or3b_1
Xhold1014 total_design.core.regFile.register\[2\]\[24\] vssd1 vssd1 vccd1 vccd1 net2330
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ net238 net2242 net440 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1025 total_design.core.regFile.register\[14\]\[10\] vssd1 vssd1 vccd1 vccd1 net2341
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 total_design.core.regFile.register\[29\]\[12\] vssd1 vssd1 vccd1 vccd1 net2352
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout286_A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1047 total_design.core.regFile.register\[13\]\[6\] vssd1 vssd1 vccd1 vccd1 net2363
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _03998_ _03999_ _01766_ vssd1 vssd1 vccd1 vccd1 total_design.core.next_instr_wait
+ sky130_fd_sc_hd__a21oi_1
Xhold1058 total_design.core.regFile.register\[13\]\[0\] vssd1 vssd1 vccd1 vccd1 net2374
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12121__B1 _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1069 total_design.core.regFile.register\[10\]\[11\] vssd1 vssd1 vccd1 vccd1 net2385
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08675_ total_design.keypad0.counter\[3\] total_design.keypad0.counter\[4\] total_design.keypad0.counter\[5\]
+ _03950_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__and4_1
XANTENNA__13742__Q total_design.core.data_bus_o\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout453_A _04117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1195_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08340__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07626_ net749 _03138_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[20\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_159_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07557_ total_design.core.regFile.register\[14\]\[19\] net862 net847 total_design.core.regFile.register\[15\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout620_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout718_A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08782__B total_design.core.data_mem.data_cpu_i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06508_ total_design.core.regFile.register\[1\]\[0\] net743 net736 net729 vssd1 vssd1
+ vccd1 vccd1 _02082_ sky130_fd_sc_hd__and4_1
XFILLER_0_91_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07488_ total_design.core.regFile.register\[30\]\[18\] net659 net624 total_design.core.regFile.register\[14\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__a22o_1
XANTENNA__07300__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09227_ _04471_ _04472_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__or2_1
XANTENNA__06654__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06439_ net971 net951 _02012_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__and3_2
XFILLER_0_133_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10309__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_X net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09158_ _04404_ _04405_ net706 vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08109_ _03600_ _03601_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__xor2_4
XFILLER_0_102_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09089_ _04234_ _04235_ net461 vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11120_ _05359_ _05378_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__xor2_2
XFILLER_0_31_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold870 total_design.core.regFile.register\[7\]\[19\] vssd1 vssd1 vccd1 vccd1 net2186
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout875_X net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold881 total_design.core.regFile.register\[10\]\[14\] vssd1 vssd1 vccd1 vccd1 net2197
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ net352 _05242_ _05305_ _05309_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__a31o_1
Xhold892 total_design.core.regFile.register\[20\]\[11\] vssd1 vssd1 vccd1 vccd1 net2208
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10044__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07906__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ net221 net2609 net417 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__mux2_1
XANTENNA__09833__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07119__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ _05803_ _05811_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__nor2_4
XANTENNA__06477__B net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10904_ _05139_ _05145_ _05142_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_28_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11884_ net897 _02188_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13623_ clknet_leaf_50_clk net1339 net1100 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10835_ total_design.core.data_bus_o\[8\] net698 vssd1 vssd1 vccd1 vccd1 _05094_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11603__S net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13554_ clknet_leaf_136_clk _01021_ net1180 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_109_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10766_ _01854_ _01857_ net930 vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09292__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10727__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14483__Q total_design.core.ctrl.instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12505_ net976 total_design.core.instr_mem.instruction_i\[16\] vssd1 vssd1 vccd1
+ vccd1 _01707_ sky130_fd_sc_hd__and2b_1
XFILLER_0_125_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10219__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13485_ clknet_leaf_6_clk _00952_ net1017 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10697_ net257 net2616 net359 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12436_ net1979 net257 net346 vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11726__A_N _05692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ net899 _03330_ _01629_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12434__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06940__B _02492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap349_A _05819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14106_ clknet_leaf_87_clk _01286_ net1248 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_11318_ _05576_ _05538_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__and2b_1
XANTENNA__07070__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12298_ net990 _04678_ net894 vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_39_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11249_ _05506_ _05507_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__or2_1
X_14037_ clknet_leaf_89_clk _01217_ net1258 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09028__B _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06790_ total_design.core.regFile.register\[4\]\[5\] net622 net572 total_design.core.regFile.register\[17\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__a22o_1
XANTENNA__12103__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08307__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11__f_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08460_ _03777_ _03783_ _03812_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_65_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07530__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07411_ net552 total_design.core.data_mem.data_cpu_i\[16\] total_design.core.ctrl.imm_32\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__a21o_1
XANTENNA_wire307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08391_ _01888_ _03747_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__and2_1
XFILLER_0_161_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_15_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_102_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07342_ total_design.core.regFile.register\[29\]\[15\] net800 net796 total_design.core.regFile.register\[11\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07273_ total_design.core.regFile.register\[7\]\[14\] net652 _02056_ total_design.core.regFile.register\[26\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__a22o_1
XANTENNA__09985__Y _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10129__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09012_ _04263_ _04264_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06224_ total_design.core.instr_mem.instruction_adr_i\[28\] total_design.core.instr_mem.instruction_adr_stored\[28\]
+ net983 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__mux2_1
XANTENNA__09918__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08747__A2_N total_design.core.data_mem.data_cpu_i\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold100 total_design.core.data_mem.data_cpu_i_reg\[13\] vssd1 vssd1 vccd1 vccd1 net1416
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06155_ net966 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__inv_2
Xhold111 total_design.core.instr_mem.instruction_adr_stored\[0\] vssd1 vssd1 vccd1
+ vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold122 total_design.core.instr_mem.instruction_adr_stored\[23\] vssd1 vssd1 vccd1
+ vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold133 total_design.core.instr_mem.instruction_adr_stored\[15\] vssd1 vssd1 vccd1
+ vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold144 total_design.core.data_mem.data_read_adr_reg2\[0\] vssd1 vssd1 vccd1 vccd1
+ net1460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 total_design.core.data_mem.data_read_adr_reg2\[2\] vssd1 vssd1 vccd1 vccd1
+ net1471 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07061__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold166 total_design.core.data_mem.data_bus_i_reg\[18\] vssd1 vssd1 vccd1 vccd1 net1482
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 total_design.core.data_mem.data_read_adr_reg2\[25\] vssd1 vssd1 vccd1 vccd1
+ net1493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold188 total_design.core.data_mem.data_cpu_i_reg\[15\] vssd1 vssd1 vccd1 vccd1 net1504
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 total_design.lcd_display.row_1\[106\] vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 net603 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_8
X_09914_ net167 net2628 net428 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__mux2_1
Xfanout613 net615 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1110_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout624 net627 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__buf_4
Xfanout635 _02061_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_4
Xfanout646 _02056_ vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09506__X _04740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ net171 net2298 net434 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__mux2_1
Xfanout657 net658 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11696__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout570_A _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 net669 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__buf_4
Xfanout679 net681 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout289_X net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ net173 total_design.core.regFile.register\[29\]\[28\] net444 vssd1 vssd1
+ vccd1 vccd1 _00099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06988_ _02537_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_126_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ total_design.key_confirm _00034_ _00032_ _03984_ vssd1 vssd1 vccd1 vccd1
+ _03986_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout456_X net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08313__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ total_design.lcd_display.cnt_500hz\[9\] _03939_ vssd1 vssd1 vccd1 vccd1 _03941_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_1_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07609_ _03119_ _03120_ _03121_ _03122_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__or4_1
XANTENNA__06875__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ _03884_ net880 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[10\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11423__S net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10620_ net179 total_design.core.regFile.register\[4\]\[27\] net367 vssd1 vssd1 vccd1
+ vccd1 _00898_ sky130_fd_sc_hd__mux2_1
X_14530__1302 vssd1 vssd1 vccd1 vccd1 net1302 _14530__1302/LO sky130_fd_sc_hd__conb_1
XFILLER_0_92_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10959__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10551_ net190 net1906 net375 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__mux2_1
XANTENNA__06627__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10039__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09828__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13270_ clknet_leaf_156_clk _00737_ net1140 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10482_ net201 net2438 net378 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__mux2_1
XANTENNA__09026__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12221_ _06067_ total_design.core.math.pc_val\[8\] net526 vssd1 vssd1 vccd1 vccd1
+ _01478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07588__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ total_design.lcd_display.row_2\[31\] _05832_ _05852_ total_design.lcd_display.row_2\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06252__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11378__B _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07052__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ total_design.core.data_bus_o\[11\] net511 _05049_ _05361_ vssd1 vssd1 vccd1
+ vccd1 _05362_ sky130_fd_sc_hd__o31a_1
XFILLER_0_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12083_ total_design.lcd_display.row_2\[60\] net348 _05847_ total_design.lcd_display.row_2\[36\]
+ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11034_ _05287_ _05288_ _05289_ _05292_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10502__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12985_ clknet_leaf_195_clk _00452_ net1010 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08304__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11936_ _05742_ _05732_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_59_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06866__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11867_ _01723_ _05723_ total_design.lcd_display.currentState\[5\] vssd1 vssd1 vccd1
+ vccd1 _05750_ sky130_fd_sc_hd__a21oi_1
X_13606_ clknet_leaf_58_clk net1331 net1125 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07768__A_N _03273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10818_ net34 total_design.core.data_bus_o\[9\] _05028_ vssd1 vssd1 vccd1 vccd1 _05077_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_138_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11798_ _03909_ _05701_ net713 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13537_ clknet_leaf_122_clk _01004_ net1169 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_10749_ net2235 net355 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07291__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13468_ clknet_leaf_28_clk _00935_ net1075 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12419_ _01674_ _01675_ net993 vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06670__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13399_ clknet_leaf_162_clk _00866_ net1166 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06251__B1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07960_ total_design.core.regFile.register\[0\]\[27\] net684 _03454_ _03458_ vssd1
+ vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__o22a_4
Xclkbuf_leaf_4_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06911_ total_design.core.regFile.register\[22\]\[7\] net677 net620 total_design.core.regFile.register\[4\]\[7\]
+ _02450_ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07891_ _03386_ _03388_ _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_147_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09630_ _04196_ _04850_ _04855_ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__o31a_1
X_06842_ _02348_ _02393_ _02391_ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__a21o_1
XANTENNA__10412__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07751__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06773_ _02334_ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09561_ _04247_ _04250_ net467 vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_104_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08512_ net933 total_design.keypad0.key_out\[10\] total_design.keypad0.key_out\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06548__D net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09492_ _03138_ net703 _04725_ net534 vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_19_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07503__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08443_ total_design.keypad0.key_out\[5\] total_design.keypad0.key_out\[4\] total_design.keypad0.key_out\[7\]
+ total_design.keypad0.key_out\[6\] vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_121_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06857__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout151_A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08374_ _03730_ _03731_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07325_ total_design.core.regFile.register\[25\]\[15\] net649 net568 total_design.core.regFile.register\[12\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__a22o_1
XANTENNA__06609__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout416_A _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1158_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07256_ _02770_ _02789_ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__nor2_1
XANTENNA__07282__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06207_ net998 net997 total_design.core.data_adr_o\[9\] vssd1 vssd1 vccd1 vccd1 _01786_
+ sky130_fd_sc_hd__o21bai_1
XANTENNA__09559__A1 _03273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07187_ total_design.core.regFile.register\[18\]\[12\] net857 _02724_ _02725_ vssd1
+ vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__a211o_1
XANTENNA__07034__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout785_A _01986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout410 net413 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__buf_6
XANTENNA__08788__A _02666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout421 _04981_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_6
Xfanout432 net433 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__buf_4
Xfanout443 _04969_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_4
Xfanout454 _04117_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11418__S net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 net466 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_2
Xfanout476 net479 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10322__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09828_ net236 net2085 net435 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__mux2_1
Xfanout487 _05007_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_4
Xfanout498 _05004_ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_6
XANTENNA__07742__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09759_ net240 net2131 net443 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout838_X net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12094__A2 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12770_ clknet_leaf_127_clk _00237_ net1192 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11721_ wishbone.curr_state\[1\] net1 wishbone.curr_state\[2\] vssd1 vssd1 vccd1
+ vccd1 _05692_ sky130_fd_sc_hd__or3b_4
XFILLER_0_139_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06848__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14440_ clknet_leaf_59_clk net1764 net1127 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11652_ _05478_ _05480_ _05674_ _05675_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__or4b_1
XFILLER_0_49_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10603_ net254 net2524 net365 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14371_ clknet_leaf_199_clk _01512_ net1001 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11583_ _05650_ net1814 net143 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13322_ clknet_leaf_21_clk _00789_ net1051 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10534_ net267 net1939 net374 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__mux2_1
XANTENNA__07273__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10465_ net282 net2107 net377 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__mux2_1
X_13253_ clknet_leaf_116_clk _00720_ net1203 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06490__B net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12204_ total_design.core.math.pc_val\[7\] total_design.core.program_count.imm_val_reg\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07025__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13184_ clknet_leaf_1_clk _00651_ net1005 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10396_ net244 net2837 net385 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__mux2_1
XANTENNA__06233__A0 total_design.core.instr_mem.instruction_adr_i\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12135_ total_design.lcd_display.row_2\[87\] _05818_ _05826_ total_design.lcd_display.row_1\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__a22o_1
XANTENNA__07981__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12066_ total_design.lcd_display.row_1\[59\] _05839_ _05848_ total_design.lcd_display.row_2\[123\]
+ _05924_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_53_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10740__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13468__RESET_B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11017_ _05247_ _05255_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__nand2_1
XANTENNA__10232__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07733__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06368__D net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12085__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12968_ clknet_leaf_172_clk _00435_ net1056 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09322__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ _03908_ _05774_ _05789_ _05794_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__a211o_1
X_12899_ clknet_leaf_8_clk _00366_ net1018 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07110_ total_design.core.regFile.register\[26\]\[11\] _02056_ net623 total_design.core.regFile.register\[4\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__a22o_1
X_08090_ total_design.core.regFile.register\[29\]\[30\] net657 net642 total_design.core.regFile.register\[19\]\[30\]
+ _03582_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload20 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_2
X_07041_ _02585_ _02586_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__and2_2
XFILLER_0_28_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload31 clknet_leaf_185_clk vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__inv_8
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10407__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload42 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__clkinv_4
Xclkload53 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__inv_16
XFILLER_0_140_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload64 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_77_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload75 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__inv_8
Xclkload86 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_100_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload97 clknet_leaf_151_clk vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_149_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11586__X _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08764__A2 _03322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08992_ net318 _04231_ _04236_ _04244_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06775__A1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07972__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07943_ total_design.core.regFile.register\[31\]\[27\] net602 net578 total_design.core.regFile.register\[27\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout199_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10142__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ total_design.core.regFile.register\[18\]\[26\] net859 net851 total_design.core.regFile.register\[9\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_3_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09931__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09613_ total_design.core.data_cpu_o\[25\] net755 _04837_ _04841_ vssd1 vssd1 vccd1
+ vccd1 _04842_ sky130_fd_sc_hd__a211o_2
XANTENNA__06559__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07017__A _02564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06825_ total_design.core.regFile.register\[26\]\[5\] net871 _02383_ _02384_ vssd1
+ vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout366_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09544_ _04765_ _04773_ _04775_ net451 vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__a31o_1
XANTENNA__12076__A2 _05840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06756_ total_design.core.regFile.register\[25\]\[4\] net647 net601 total_design.core.regFile.register\[31\]\[4\]
+ _02316_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13750__Q total_design.core.data_bus_o\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06687_ total_design.core.regFile.register\[30\]\[3\] net838 _02243_ _01932_ vssd1
+ vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09475_ _04709_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout154_X net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout533_A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08426_ total_design.keypad0.key_out\[11\] total_design.keypad0.key_out\[8\] vssd1
+ vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08357_ total_design.keypad0.key_out\[1\] total_design.keypad0.key_out\[2\] total_design.keypad0.key_out\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08790__B _02868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_33_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07308_ _02818_ _02838_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__and2b_1
X_08288_ net1492 net941 _03678_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[1\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_172_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1550_A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10317__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07239_ total_design.core.regFile.register\[23\]\[13\] net813 net805 total_design.core.regFile.register\[8\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12536__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10250_ net205 net2459 net500 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__mux2_1
XANTENNA__07007__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08755__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ net183 net2382 net395 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1205 net1206 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__clkbuf_4
Xfanout1216 net1219 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__clkbuf_4
Xfanout1227 net1232 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout955_X net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1238 net1239 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__clkbuf_4
Xfanout240 net243 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_2
Xfanout1249 net1251 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__clkbuf_4
Xfanout251 net252 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout262 net264 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_2
X_13940_ clknet_leaf_98_clk _01120_ net1244 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[86\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout273 net274 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11375__C _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11511__A1 _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout284 net287 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_2
Xfanout295 net297 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_2
XANTENNA__09841__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06469__C net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ clknet_leaf_68_clk total_design.core.ctrl.imm_32\[10\] net1111 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08965__B _02917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12822_ clknet_leaf_153_clk _00289_ net1136 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10559__Y _05013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12753_ clknet_leaf_151_clk _00220_ net1145 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08140__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06485__B net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11704_ net8 net934 net877 net1824 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__o22a_1
XANTENNA__07494__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12684_ clknet_leaf_166_clk _00151_ net1157 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14423_ clknet_leaf_34_clk total_design.core.data_out_INSTR\[18\] net1067 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[18\] sky130_fd_sc_hd__dfrtp_1
X_11635_ _05680_ net1688 net136 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11611__S net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14354_ clknet_leaf_45_clk _00023_ net1086 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07246__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11566_ _05632_ net1848 net144 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10735__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14491__Q total_design.core.ctrl.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13305_ clknet_leaf_197_clk _00772_ net1007 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10517_ net195 net2043 net480 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14285_ net987 _01461_ net1082 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11497_ net1572 _05665_ net149 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13236_ clknet_leaf_142_clk _00703_ net1176 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10448_ net208 net2152 net381 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08746__A2 _03178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ clknet_leaf_161_clk _00634_ net1153 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12442__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10379_ net213 total_design.core.regFile.register\[11\]\[17\] net484 vssd1 vssd1
+ vccd1 vccd1 _00664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07954__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11750__B2 total_design.core.data_bus_o\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12118_ total_design.lcd_display.row_2\[94\] _05837_ _05846_ total_design.lcd_display.row_2\[102\]
+ _05973_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_72_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13098_ clknet_leaf_22_clk _00565_ net1049 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12049_ net124 net709 _05894_ _05908_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__o22a_1
XANTENNA__11502__A1 _05655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07706__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09751__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__B _02818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06610_ _02170_ _02171_ _02172_ _02173_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__or4_1
X_07590_ total_design.core.regFile.register\[2\]\[20\] net636 net569 total_design.core.regFile.register\[17\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12058__A2 _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09459__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07124__X _02666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06541_ _02106_ net469 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__nand2_1
XANTENNA__08594__C net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06395__B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06472_ net741 net728 net726 vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__and3_1
X_09260_ _04503_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__inv_2
XANTENNA__07485__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09707__A_N net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ _03664_ _03665_ _03667_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__or3_1
XANTENNA__06693__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09191_ net461 _04389_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10926__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11521__S net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08142_ total_design.core.regFile.register\[9\]\[31\] net664 net621 total_design.core.regFile.register\[4\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__a22o_1
XANTENNA__07237__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08073_ total_design.core.regFile.register\[25\]\[30\] net844 net833 total_design.core.regFile.register\[31\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__a22o_1
Xclkload120 clknet_leaf_170_clk vssd1 vssd1 vccd1 vccd1 clkload120/Y sky130_fd_sc_hd__inv_8
XFILLER_0_153_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload131 clknet_leaf_149_clk vssd1 vssd1 vccd1 vccd1 clkload131/Y sky130_fd_sc_hd__inv_8
XANTENNA__10137__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload142 clknet_leaf_135_clk vssd1 vssd1 vccd1 vccd1 clkload142/Y sky130_fd_sc_hd__clkinv_2
Xclkload153 clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 clkload153/Y sky130_fd_sc_hd__inv_8
X_07024_ total_design.core.regFile.register\[10\]\[9\] net836 net825 total_design.core.regFile.register\[19\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a22o_1
XANTENNA__06561__D net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09926__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload164 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 clkload164/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_168_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload175 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 clkload175/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_168_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07945__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13745__Q total_design.core.data_bus_o\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ net336 _02613_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__or2_1
XANTENNA__08131__A _03622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 total_design.core.data_mem.data_read_adr_reg\[10\] vssd1 vssd1 vccd1 vccd1
+ net1331 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout483_A _05011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold26 total_design.core.data_mem.data_read_adr_reg\[28\] vssd1 vssd1 vccd1 vccd1
+ net1342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 total_design.core.data_mem.data_bus_i_reg\[2\] vssd1 vssd1 vccd1 vccd1 net1353
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ total_design.core.regFile.register\[1\]\[27\] net828 net780 total_design.core.regFile.register\[27\]\[27\]
+ _03425_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__a221o_1
Xhold48 total_design.core.data_mem.data_cpu_i_reg\[12\] vssd1 vssd1 vccd1 vccd1 net1364
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 total_design.core.math.pc_val\[10\] vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ total_design.core.regFile.register\[19\]\[25\] net641 net618 total_design.core.regFile.register\[10\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__B total_design.core.data_mem.data_cpu_i\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11800__B1_N net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06808_ total_design.core.regFile.register\[11\]\[5\] net796 net769 total_design.core.regFile.register\[7\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__a22o_1
XANTENNA__10600__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12049__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07788_ total_design.core.regFile.register\[26\]\[24\] net870 net862 total_design.core.regFile.register\[14\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12954__RESET_B net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09527_ net507 _04759_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06739_ _02296_ _02298_ _02300_ _02302_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08122__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_X net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07476__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09458_ _04507_ _04687_ _04693_ net289 _04689_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__o221a_1
XFILLER_0_54_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08409_ _03762_ _03763_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__xor2_1
XANTENNA__06684__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10836__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09389_ _02892_ net508 net446 _02891_ _04627_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__o221a_1
XANTENNA__11431__S net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11420_ net1756 _05618_ net157 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07228__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07210__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11351_ net510 net304 vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__or2_2
XFILLER_0_132_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10047__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08976__A2 _02564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09836__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10302_ net275 net2363 net494 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__mux2_1
X_14070_ clknet_leaf_100_clk _01250_ net1237 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_89_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11282_ _05481_ _05494_ _05495_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__nand3_2
XFILLER_0_132_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08189__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ clknet_leaf_20_clk _00488_ net1026 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10233_ net268 net2641 net501 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__mux2_1
XANTENNA__12115__X _05971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06260__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1002 net1006 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_2
X_10164_ net251 net2063 net396 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__mux2_1
Xfanout1013 net1014 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07400__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1024 net1027 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_4
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1046 net1051 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_4
Xfanout1057 net1058 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__clkbuf_4
X_10095_ net261 total_design.core.regFile.register\[19\]\[8\] net404 vssd1 vssd1 vccd1
+ vccd1 _00399_ sky130_fd_sc_hd__mux2_1
Xfanout1068 net1069 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1079 net1080 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__clkbuf_2
X_13923_ clknet_leaf_88_clk _01103_ net1260 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11606__S net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13854_ clknet_leaf_54_clk _01062_ net1117 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10510__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12805_ clknet_leaf_117_clk _00272_ net1212 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14486__Q total_design.core.ctrl.instruction\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13785_ clknet_leaf_56_clk total_design.core.data_mem.stored_data_adr\[28\] net1114
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10997_ _05250_ _05255_ _05247_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__a21o_1
XANTENNA__08113__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12736_ clknet_leaf_193_clk _00203_ net1012 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06675__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ clknet_leaf_146_clk _00134_ net1177 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12437__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14406_ clknet_leaf_38_clk total_design.core.data_out_INSTR\[1\] net1078 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[1\] sky130_fd_sc_hd__dfrtp_1
X_11618_ _05630_ net1634 net140 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07219__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09613__B1 _04837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12598_ clknet_leaf_156_clk _00065_ net1142 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14337_ clknet_leaf_54_clk _01498_ net1110 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[28\]
+ sky130_fd_sc_hd__dfstp_1
X_11549_ net1551 _05633_ net147 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold507 net40 vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 total_design.keypad0.key_clk vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06381__D net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold529 total_design.core.math.pc_val\[6\] vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14268_ clknet_leaf_46_clk _00000_ net1088 vssd1 vssd1 vccd1 vccd1 wishbone.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_123_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmax_cap248 _05547_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_1
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ clknet_leaf_7_clk _00686_ net1016 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14199_ clknet_leaf_80_clk _01379_ net1221 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07927__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 total_design.core.regFile.register\[3\]\[9\] vssd1 vssd1 vccd1 vccd1 net2523
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ _04010_ _04011_ _04012_ _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__or4_1
Xhold1218 total_design.core.regFile.register\[1\]\[16\] vssd1 vssd1 vccd1 vccd1 net2534
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 total_design.core.regFile.register\[27\]\[31\] vssd1 vssd1 vccd1 vccd1 net2545
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07711_ total_design.core.regFile.register\[23\]\[22\] net679 net617 total_design.core.regFile.register\[10\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__a22o_1
X_08691_ total_design.keypad0.counter\[13\] _03956_ net2015 vssd1 vssd1 vccd1 vccd1
+ _03964_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_201_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_201_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07642_ total_design.core.regFile.register\[26\]\[21\] net870 net843 total_design.core.regFile.register\[25\]\[21\]
+ _03153_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__a221o_1
XANTENNA__10420__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07573_ _03044_ _03088_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__xor2_4
XANTENNA__08104__B1 total_design.core.ctrl.imm_32\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09312_ net313 _04356_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__nand2_1
XANTENNA__14200__RESET_B net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06556__D net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06524_ total_design.core.regFile.register\[17\]\[0\] net570 _02093_ _02079_ _02082_
+ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07458__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ net318 _04231_ _04487_ net297 vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__a211o_1
XFILLER_0_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06455_ _01924_ _02020_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_157_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09174_ net298 _04410_ _04420_ _04421_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__o211a_1
X_06386_ total_design.core.regFile.register\[1\]\[0\] net922 net949 net910 vssd1 vssd1
+ vccd1 vccd1 _01962_ sky130_fd_sc_hd__and4_1
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08125_ total_design.core.regFile.register\[26\]\[31\] net870 net768 total_design.core.regFile.register\[7\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07615__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07965__A _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ total_design.core.regFile.register\[0\]\[29\] net682 _03546_ _03550_ vssd1
+ vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07630__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout698_A net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07007_ total_design.core.regFile.register\[26\]\[9\] net646 net635 total_design.core.regFile.register\[16\]\[9\]
+ _02554_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1026_X net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_X net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_A _01941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ net469 _02182_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__nor2_1
X_07909_ total_design.core.regFile.register\[27\]\[26\] net578 _03408_ _03409_ vssd1
+ vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__a211o_1
XANTENNA__07146__A1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout653_X net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08889_ net334 net311 vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__and2_1
XANTENNA__11426__S net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ _05157_ _05159_ _05161_ _05167_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__a31o_1
XANTENNA__10330__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10851_ _05108_ _05109_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout820_X net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11372__D _05630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13570_ clknet_leaf_41_clk total_design.core.data_mem.data_bus_i\[6\] net1090 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_160_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07449__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10782_ total_design.core.data_bus_o\[17\] total_design.core.data_bus_o\[24\] total_design.core.data_bus_o\[26\]
+ total_design.core.data_bus_o\[27\] net696 vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__o41a_1
XFILLER_0_13_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11650__A0 _05651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06657__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12521_ net974 total_design.core.instr_mem.instruction_i\[24\] vssd1 vssd1 vccd1
+ vccd1 _01715_ sky130_fd_sc_hd__and2b_1
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12452_ net2778 net202 net345 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11403_ _05380_ net304 vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_175_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12383_ _01641_ _01642_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__or2_1
X_14122_ clknet_leaf_86_clk _01302_ net1247 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11334_ _05591_ _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07082__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14053_ clknet_leaf_92_clk _01233_ net1262 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11265_ _05434_ _05436_ _05522_ _05523_ _05431_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10505__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ clknet_leaf_167_clk _00471_ net1156 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10216_ _04804_ net2868 net389 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__mux2_1
XANTENNA__09374__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11196_ _05449_ _05451_ _05453_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__nand3_2
XANTENNA__06188__A2 net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10147_ net182 net1942 net400 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10078_ net190 net2283 net407 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12805__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13906_ clknet_leaf_87_clk _01086_ net1250 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10240__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09314__B net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07688__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13837_ clknet_leaf_58_clk _01045_ net1126 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06896__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_128_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06376__D net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13768_ clknet_leaf_59_clk total_design.core.data_mem.stored_data_adr\[11\] net1126
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11641__A0 _05609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06648__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12719_ clknet_leaf_146_clk _00186_ net1152 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_13699_ clknet_leaf_40_clk total_design.core.data_mem.stored_read_data\[6\] net1090
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06240_ net998 net997 total_design.core.data_adr_o\[31\] vssd1 vssd1 vccd1 vccd1
+ _01819_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_135_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07860__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09598__C1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06171_ total_design.core.data_cpu_o\[6\] vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold304 total_design.lcd_display.row_1\[2\] vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07073__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold315 total_design.core.math.pc_val\[5\] vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07612__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold326 total_design.lcd_display.row_1\[52\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold337 net74 vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold348 total_design.lcd_display.row_2\[107\] vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06820__B1 _01969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09930_ net236 net2426 net422 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__mux2_1
Xhold359 total_design.lcd_display.row_2\[85\] vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10415__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09048__Y _04300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11100__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout806 net809 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_8
Xfanout817 net818 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_4
X_09861_ net241 net2516 net430 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout828 net830 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__buf_4
Xfanout839 net841 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__buf_4
X_08812_ _02367_ _02388_ _04066_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__a21o_1
X_09792_ net241 net2224 net441 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__mux2_1
Xhold1004 total_design.core.regFile.register\[7\]\[9\] vssd1 vssd1 vccd1 vccd1 net2320
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1015 total_design.core.regFile.register\[21\]\[12\] vssd1 vssd1 vccd1 vccd1 net2331
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1026 total_design.core.regFile.register\[22\]\[2\] vssd1 vssd1 vccd1 vccd1 net2342
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ _02025_ _03467_ total_design.core.data_mem.data_write_adr_i\[11\] vssd1 vssd1
+ vccd1 vccd1 _03999_ sky130_fd_sc_hd__o21ba_1
Xhold1037 total_design.core.regFile.register\[11\]\[8\] vssd1 vssd1 vccd1 vccd1 net2353
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 total_design.core.regFile.register\[11\]\[12\] vssd1 vssd1 vccd1 vccd1 net2364
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 total_design.core.regFile.register\[12\]\[21\] vssd1 vssd1 vccd1 vccd1 net2375
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout181_A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_A _04315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10150__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08674_ total_design.keypad0.counter\[3\] _03950_ vssd1 vssd1 vccd1 vccd1 _03951_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07679__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07625_ _03093_ _03136_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout446_A _04189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07556_ total_design.core.regFile.register\[30\]\[19\] net839 _03072_ _03073_ vssd1
+ vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__a211o_1
XANTENNA__11632__A0 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06507_ net742 net736 net728 vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07487_ _03001_ _03003_ _03005_ _03007_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout613_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout234_X net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09226_ total_design.core.math.pc_val\[8\] _04448_ vssd1 vssd1 vccd1 vccd1 _04472_
+ sky130_fd_sc_hd__nor2_1
X_06438_ total_design.core.ctrl.instruction\[4\] net973 net972 vssd1 vssd1 vccd1 vccd1
+ _02013_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_1_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07851__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09157_ _02390_ _04403_ _02441_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06369_ net926 net948 net916 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07064__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08108_ _03507_ _03510_ _03555_ _03553_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__o31a_2
XFILLER_0_82_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07603__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09088_ net463 _04239_ _04338_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_169_Right_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout982_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08039_ total_design.core.regFile.register\[7\]\[29\] net651 net644 total_design.core.regFile.register\[26\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__a22o_1
XANTENNA__10325__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold860 total_design.core.regFile.register\[3\]\[16\] vssd1 vssd1 vccd1 vccd1 net2176
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold871 total_design.core.regFile.register\[3\]\[28\] vssd1 vssd1 vccd1 vccd1 net2187
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 total_design.core.regFile.register\[13\]\[9\] vssd1 vssd1 vccd1 vccd1 net2198
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11050_ _05033_ _05046_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__nor2_1
Xhold893 total_design.core.regFile.register\[12\]\[31\] vssd1 vssd1 vccd1 vccd1 net2209
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_X net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ net224 net2274 net416 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14193__RESET_B net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09513__C1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1560 net87 vssd1 vssd1 vccd1 vccd1 net2876 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10060__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11952_ _05809_ _05813_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06477__C net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10903_ _05139_ _05145_ _05142_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__or3b_1
XANTENNA__06878__B1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ total_design.core.math.pc_val\[0\] _05763_ _05759_ vssd1 vssd1 vccd1 vccd1
+ _01444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08973__B _02718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13622_ clknet_leaf_50_clk net1333 net1100 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10834_ _05076_ _05079_ _05085_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__and3_1
XANTENNA__09816__A0 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06774__A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11623__A0 _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13553_ clknet_leaf_148_clk _01020_ net1146 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10765_ _01887_ _05023_ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__nor2_1
XANTENNA__08095__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06493__B _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12504_ net974 total_design.core.ctrl.instruction\[15\] net881 _01706_ vssd1 vssd1
+ vccd1 vccd1 _01554_ sky130_fd_sc_hd__a22o_1
XANTENNA__07842__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13484_ clknet_leaf_168_clk _00951_ net1158 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10696_ net280 total_design.core.regFile.register\[1\]\[4\] net357 vssd1 vssd1 vccd1
+ vccd1 _00971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12435_ net2025 net281 net344 vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07055__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12366_ net991 _04819_ _01628_ net894 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_130_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10743__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14105_ clknet_leaf_96_clk _01285_ net1257 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_11317_ _05571_ _05573_ _05575_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06802__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10235__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12297_ _06132_ _06133_ _06131_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__o21ai_1
X_14036_ clknet_leaf_99_clk _01216_ net1229 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[118\]
+ sky130_fd_sc_hd__dfrtp_1
X_11248_ _05408_ _05498_ _05504_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__and3_1
XANTENNA__09062__A2_N net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12450__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ _05434_ _05436_ _05431_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08307__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06869__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08883__B _02666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07410_ total_design.core.regFile.register\[0\]\[16\] net876 _02920_ _02936_ vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[16\] sky130_fd_sc_hd__o22a_4
X_08390_ _01732_ _03719_ _03744_ _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_174_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11614__A0 _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07341_ total_design.core.regFile.register\[24\]\[15\] net792 _02870_ vssd1 vssd1
+ vccd1 vccd1 _02871_ sky130_fd_sc_hd__a21o_1
XANTENNA__08086__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07272_ total_design.core.regFile.register\[23\]\[14\] net678 net589 total_design.core.regFile.register\[1\]\[14\]
+ _02800_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__a221o_1
XANTENNA__07833__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09011_ net472 net306 vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06223_ total_design.core.data_adr_o\[14\] _01801_ net963 vssd1 vssd1 vccd1 vccd1
+ _01802_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_171_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10493__X _05011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06154_ total_design.core.ctrl.instruction\[21\] vssd1 vssd1 vccd1 vccd1 _01737_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_124_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold101 total_design.core.data_mem.data_cpu_i_reg\[1\] vssd1 vssd1 vccd1 vccd1 net1417
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 total_design.core.data_mem.data_bus_i_reg\[31\] vssd1 vssd1 vccd1 vccd1 net1428
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 total_design.core.data_mem.data_bus_i_reg\[25\] vssd1 vssd1 vccd1 vccd1 net1439
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 total_design.core.data_mem.data_bus_i_reg\[17\] vssd1 vssd1 vccd1 vccd1 net1450
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 total_design.core.data_mem.data_bus_i_reg\[12\] vssd1 vssd1 vccd1 vccd1 net1461
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10145__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold156 total_design.core.data_mem.data_read_adr_reg2\[7\] vssd1 vssd1 vccd1 vccd1
+ net1472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 total_design.core.data_mem.data_bus_i_reg\[27\] vssd1 vssd1 vccd1 vccd1 net1483
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 total_design.core.data_mem.data_read_adr_reg2\[17\] vssd1 vssd1 vccd1 vccd1
+ net1494 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ net170 net2620 net426 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__mux2_1
XANTENNA__09934__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09338__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold189 net54 vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _02076_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout614 net615 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_4
XANTENNA_fanout396_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout625 net627 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 net639 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09743__C1 _04963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09844_ net173 net2832 net437 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__mux2_1
Xfanout647 net650 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_8
Xfanout658 _02052_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_4
Xfanout669 _02046_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__buf_4
X_09775_ net178 net2099 net445 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__mux2_1
X_06987_ _02515_ _02535_ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__and2b_1
XANTENNA__13753__Q total_design.core.data_bus_o\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout563_A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06578__B net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout184_X net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06572__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08657_ total_design.lcd_display.cnt_500hz\[9\] _03939_ vssd1 vssd1 vccd1 vccd1 _03940_
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout730_A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout828_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08793__B _02718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07608_ total_design.core.regFile.register\[11\]\[20\] net794 net759 total_design.core.regFile.register\[21\]\[20\]
+ _03113_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08588_ _03873_ net880 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[9\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11605__A0 _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07539_ total_design.core.regFile.register\[9\]\[19\] net664 net567 total_design.core.regFile.register\[12\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__a22o_1
XANTENNA__08077__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10959__A2 _05184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_10__f_clk_X clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ net194 net2784 net373 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06881__X total_design.core.data_mem.data_cpu_i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09209_ _02539_ _04454_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07696__Y _03206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10481_ net206 net2863 net377 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12220_ net898 _02540_ _06065_ _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__o22a_1
XANTENNA__07037__B1 total_design.core.ctrl.imm_32\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout985_X net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ total_design.lcd_display.row_2\[111\] _05834_ _05849_ total_design.lcd_display.row_2\[55\]
+ _06005_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__a221o_1
XANTENNA__10055__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11378__C _05636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06796__C1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11102_ _01871_ _01883_ _05059_ _01900_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__or4b_2
XANTENNA__09844__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12082_ total_design.lcd_display.row_1\[44\] _05821_ _05826_ total_design.lcd_display.row_1\[20\]
+ _05939_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__a221o_1
XANTENNA__14374__RESET_B net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold690 total_design.core.regFile.register\[22\]\[14\] vssd1 vssd1 vccd1 vccd1 net2006
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08968__B _02770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ net350 _05291_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__nor2_1
XANTENNA__08001__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06488__B net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12097__B1 _05840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12984_ clknet_leaf_138_clk _00451_ net1184 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1390 total_design.core.regFile.register\[23\]\[16\] vssd1 vssd1 vccd1 vccd1 net2706
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11935_ total_design.keypad0.key_out\[15\] net529 net475 total_design.keypad0.key_out\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__a22o_1
XANTENNA__11614__S net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11866_ total_design.lcd_display.currentState\[3\] _05749_ net709 vssd1 vssd1 vccd1
+ vccd1 _01441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10738__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13605_ clknet_leaf_62_clk net1321 net1125 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10817_ _05068_ _05075_ _05072_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08068__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11797_ total_design.lcd_display.cnt_20ms\[0\] total_design.lcd_display.cnt_20ms\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13536_ clknet_leaf_192_clk _01003_ net1033 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07276__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07815__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10748_ total_design.core.regFile.register\[0\]\[23\] net353 vssd1 vssd1 vccd1 vccd1
+ _01022_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13467_ clknet_leaf_150_clk _00934_ net1148 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12445__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10679_ net207 net2225 net361 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12021__B1 _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11882__A1_N net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12418_ total_design.core.math.pc_val\[29\] net989 _01668_ vssd1 vssd1 vccd1 vccd1
+ _01675_ sky130_fd_sc_hd__a21bo_1
X_13398_ clknet_leaf_153_clk _00865_ net1138 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12349_ _01604_ _01608_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09754__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08878__B _02718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14019_ clknet_leaf_90_clk _01199_ net1260 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[101\]
+ sky130_fd_sc_hd__dfrtp_1
X_06910_ total_design.core.regFile.register\[21\]\[7\] net600 _02463_ net689 vssd1
+ vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__a211o_1
X_07890_ total_design.core.regFile.register\[11\]\[26\] net795 _03389_ _03391_ vssd1
+ vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_147_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08597__C net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06841_ total_design.core.ctrl.instruction\[18\] net887 _02149_ _02398_ _02397_ vssd1
+ vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[6\] sky130_fd_sc_hd__a221o_2
XANTENNA__06398__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12088__B1 _05829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09560_ _03279_ net509 net448 _03278_ _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__o221a_1
X_06772_ total_design.core.regFile.register\[0\]\[4\] net682 _02329_ _02333_ vssd1
+ vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_104_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08511_ _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__inv_2
X_09491_ net703 _04724_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_19_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11524__S net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08442_ _03710_ _03796_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[5\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_121_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08373_ _03725_ _03729_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_173_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09929__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07267__B1 _02076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06564__D net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07324_ total_design.core.regFile.register\[23\]\[15\] net680 net617 total_design.core.regFile.register\[10\]\[15\]
+ _02852_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07806__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07255_ _02789_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06206_ _01782_ _01784_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_30_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07019__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12012__B1 _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07186_ total_design.core.regFile.register\[25\]\[12\] net842 net830 total_design.core.regFile.register\[1\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__a22o_1
XANTENNA__13748__Q total_design.core.data_bus_o\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1220_A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10574__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06242__A1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09664__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout680_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 _04990_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_6
Xfanout411 net413 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_6
XANTENNA__08788__B net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07990__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06793__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout399_X net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 net425 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_6
XANTENNA_fanout778_A _01990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10603__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout433 _04975_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_8
Xfanout444 _04969_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_6
Xfanout455 _04117_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_8
Xfanout466 _02184_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_2
Xfanout477 net478 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_6
X_09827_ net243 net2327 net435 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__mux2_1
Xfanout488 net491 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_6
XANTENNA_fanout945_A _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout566_X net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout499 _05004_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_4
XANTENNA__12079__B1 _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ net253 net2572 net442 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__mux2_1
X_08709_ _00020_ total_design.keypad0.counter\[1\] _03972_ _03973_ vssd1 vssd1 vccd1
+ vccd1 _03974_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_61_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ _03556_ _04892_ _04913_ net707 vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__o211a_1
XANTENNA__11434__S net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11720_ net26 net934 net877 net2634 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07213__A total_design.core.ctrl.instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11651_ _05630_ net1616 net135 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout900_X net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09247__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11054__A1 total_design.core.data_bus_o\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09839__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10602_ net251 net2637 net367 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__mux2_1
X_14370_ clknet_leaf_117_clk _01511_ net1161 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11582_ _05633_ net1815 net144 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13321_ clknet_leaf_4_clk _00788_ net1023 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10533_ net273 net2763 net376 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_9__f_clk_X clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12003__B1 _05848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13252_ clknet_leaf_105_clk _00719_ net1233 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06263__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ net268 net2124 net378 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12203_ total_design.core.math.pc_val\[7\] total_design.core.program_count.imm_val_reg\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__nand2_1
XANTENNA__12649__RESET_B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13183_ clknet_leaf_154_clk _00650_ net1136 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10395_ net284 net2698 net385 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__mux2_1
XANTENNA__06769__C1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12134_ _05974_ _05976_ _05989_ net709 net2815 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_36_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07430__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09427__X _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11609__S net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12065_ total_design.lcd_display.row_2\[107\] _05834_ _05850_ total_design.lcd_display.row_2\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__a22o_1
XANTENNA__10513__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11016_ net520 _05271_ _05273_ _05269_ _05270_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__a32o_1
XANTENNA__14489__Q total_design.core.ctrl.instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06786__X _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09162__X _04410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ clknet_leaf_177_clk _00434_ net1047 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11918_ net1000 _05791_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__nor2_1
XANTENNA__07497__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09322__B _04563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12490__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12898_ clknet_leaf_126_clk _00365_ net1192 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11849_ total_design.lcd_display.currentState\[3\] _05734_ vssd1 vssd1 vccd1 vccd1
+ _05735_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07249__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06384__D net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07410__X total_design.core.data_mem.data_cpu_i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_109_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13519_ clknet_leaf_160_clk _00986_ net1151 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14499_ clknet_leaf_36_clk _01566_ net1071 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[27\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkload10 clknet_leaf_194_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_8
XFILLER_0_70_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07040_ _02586_ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload21 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__clkinv_2
Xclkload32 clknet_leaf_186_clk vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload43 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__inv_8
XFILLER_0_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload54 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload65 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload76 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_51_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload87 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_140_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload98 clknet_leaf_152_clk vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__07421__B1 total_design.core.ctrl.instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08991_ net326 _04243_ net318 vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06775__A2 total_design.core.data_mem.data_cpu_i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11519__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07942_ total_design.core.regFile.register\[19\]\[27\] net642 net609 total_design.core.regFile.register\[18\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__a22o_1
XANTENNA__10423__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07873_ net749 _03375_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[25\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_173_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09612_ net903 _04840_ _02750_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_3_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06824_ total_design.core.regFile.register\[24\]\[5\] net792 net781 total_design.core.regFile.register\[27\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_123_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06559__D net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09543_ _03227_ _04189_ _04774_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__o21a_1
X_06755_ total_design.core.regFile.register\[7\]\[4\] net651 net608 total_design.core.regFile.register\[18\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__a22o_1
XANTENNA__09477__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout261_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_A _05017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07488__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ _04668_ _04708_ net468 vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__mux2_1
X_06686_ total_design.core.regFile.register\[11\]\[3\] net795 _02251_ _02252_ vssd1
+ vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a211o_1
X_08425_ total_design.keypad0.key_out\[11\] total_design.keypad0.key_out\[8\] vssd1
+ vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout147_X net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08356_ _03714_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload4 clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__clkinv_8
X_07307_ _02838_ _02818_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08287_ total_design.core.data_mem.data_write_adr_reg\[1\] net549 net541 total_design.core.data_mem.data_read_adr_reg\[1\]
+ net945 vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__a221o_1
XANTENNA__07660__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07238_ total_design.core.regFile.register\[18\]\[13\] net857 net834 total_design.core.regFile.register\[10\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07169_ total_design.core.regFile.register\[10\]\[12\] net619 net576 total_design.core.regFile.register\[24\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10180_ net186 net2693 net395 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06766__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1206 net1211 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__clkbuf_4
Xfanout1217 net1219 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10333__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
Xfanout1228 net1231 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout241 net243 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_2
Xfanout1239 net1240 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout252 _04496_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout850_X net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout263 net264 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_31_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout274 net275 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11375__D _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout948_X net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout285 net287 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_2
Xfanout296 net297 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_2
X_13870_ clknet_leaf_68_clk total_design.core.ctrl.imm_32\[9\] net1111 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[9\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06469__D net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07191__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12821_ clknet_leaf_158_clk _00288_ net1141 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07479__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ clknet_leaf_186_clk _00219_ net1037 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06258__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06485__C net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11703_ net7 net936 net879 net1857 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__a22o_1
X_12683_ clknet_leaf_108_clk _00150_ net1224 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08981__B _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14422_ clknet_leaf_32_clk total_design.core.data_out_INSTR\[17\] net1062 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[17\] sky130_fd_sc_hd__dfrtp_1
X_11634_ _05655_ net1729 net133 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14353_ clknet_leaf_45_clk _00022_ net1086 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11565_ _05670_ net1664 net143 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__mux2_1
XANTENNA__10508__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ clknet_leaf_136_clk _00771_ net1178 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10516_ net198 net2092 net482 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14284_ net987 _01460_ net1083 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_134_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11496_ net1584 _05663_ net152 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13235_ clknet_leaf_182_clk _00702_ net1043 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10447_ net212 net2054 net382 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07403__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ clknet_leaf_189_clk _00633_ net1030 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10378_ net220 net2699 net486 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__mux2_1
XANTENNA__10751__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06757__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12117_ total_design.lcd_display.row_2\[86\] _05818_ _05832_ total_design.lcd_display.row_2\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__a22o_1
XANTENNA__11750__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10243__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13097_ clknet_leaf_192_clk _00564_ net1033 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12048_ _05898_ _05900_ _05902_ _05907_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__or4_1
XANTENNA__08903__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06379__D net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07182__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13999_ clknet_leaf_84_clk _01179_ net1245 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06676__B net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06540_ _02106_ net469 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10198__B net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06471_ _01924_ net901 _02018_ total_design.core.ctrl.instruction\[18\] total_design.core.ctrl.instruction\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__o311a_1
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08210_ total_design.core.data_mem.data_read_adr_reg\[13\] total_design.core.data_mem.data_read_adr_reg\[12\]
+ total_design.core.data_mem.data_read_adr_reg\[15\] total_design.core.data_mem.data_read_adr_reg\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__or4_1
XFILLER_0_146_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09190_ _04435_ _04436_ net318 vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10926__B _05184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08141_ total_design.core.regFile.register\[8\]\[31\] net594 net590 total_design.core.regFile.register\[1\]\[31\]
+ _03631_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10418__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07642__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08072_ total_design.core.regFile.register\[11\]\[30\] net796 net778 total_design.core.regFile.register\[22\]\[30\]
+ _03565_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__a221o_1
Xclkload110 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 clkload110/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_15_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload121 clknet_leaf_136_clk vssd1 vssd1 vccd1 vccd1 clkload121/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_116_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload132 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 clkload132/Y sky130_fd_sc_hd__inv_6
Xclkload143 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 clkload143/Y sky130_fd_sc_hd__inv_6
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload154 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 clkload154/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07023_ total_design.core.regFile.register\[3\]\[9\] net868 _02567_ _02569_ _02570_
+ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_168_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload165 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 clkload165/Y sky130_fd_sc_hd__inv_6
Xclkload176 clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 clkload176/Y sky130_fd_sc_hd__inv_8
XFILLER_0_113_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09508__A _03112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08974_ _04225_ _04226_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__nand2_1
Xhold16 total_design.core.data_mem.data_read_adr_reg\[29\] vssd1 vssd1 vccd1 vccd1
+ net1332 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09147__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold27 total_design.core.data_mem.data_read_adr_reg\[19\] vssd1 vssd1 vccd1 vccd1
+ net1343 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ total_design.core.regFile.register\[11\]\[27\] net796 net788 total_design.core.regFile.register\[13\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__a22o_1
Xhold38 total_design.core.data_mem.data_cpu_i_reg\[14\] vssd1 vssd1 vccd1 vccd1 net1354
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 total_design.core.data_mem.data_cpu_i_reg\[7\] vssd1 vssd1 vccd1 vccd1 net1365
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__A1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09698__B2 _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ total_design.core.regFile.register\[22\]\[25\] net675 net586 total_design.core.regFile.register\[28\]\[25\]
+ _03358_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__a221o_1
XANTENNA__07173__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06807_ _02351_ _02352_ _02366_ net685 total_design.core.regFile.register\[0\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__o32a_4
X_07787_ total_design.core.regFile.register\[18\]\[24\] net858 net807 total_design.core.regFile.register\[5\]\[24\]
+ _03292_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout264_X net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06920__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ _04755_ _04758_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__or2_2
X_06738_ total_design.core.regFile.register\[24\]\[4\] net790 net775 total_design.core.regFile.register\[22\]\[4\]
+ _02301_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09457_ _04597_ _04691_ net327 vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout810_A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06669_ net554 _02211_ _02235_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a21oi_1
X_08408_ _03762_ _03763_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07881__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ _02890_ net504 vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08339_ total_design.core.data_mem.data_write_adr_reg\[27\] net546 net538 total_design.core.data_mem.data_read_adr_reg\[27\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11350_ total_design.core.data_bus_o\[21\] net697 net303 _05608_ net510 vssd1 vssd1
+ vccd1 vccd1 _05609_ sky130_fd_sc_hd__a221o_4
XANTENNA__07633__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout898_X net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10301_ net258 net2001 net494 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11281_ _05498_ _05504_ _05539_ _05488_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__a31o_1
XANTENNA__10852__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13020_ clknet_leaf_28_clk _00487_ net1074 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10232_ net278 net2261 net501 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1003 net1006 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10063__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10163_ net262 net2498 net396 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__mux2_1
Xfanout1014 net1015 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09852__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1025 net1026 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_4
Xfanout1036 net1059 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input37_A gpio_in[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11954__Y _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 net1051 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__clkbuf_4
X_10094_ net267 net1947 net402 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__mux2_1
Xfanout1058 net1059 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__clkbuf_2
Xfanout1069 net1081 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13922_ clknet_leaf_87_clk _01102_ net1250 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11496__A1 _05663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13029__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06777__A _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07164__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09153__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13853_ clknet_leaf_54_clk _01061_ net1109 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06372__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06911__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06496__B net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12804_ clknet_leaf_128_clk _00271_ net1193 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13784_ clknet_leaf_50_clk total_design.core.data_mem.stored_data_adr\[27\] net1101
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[27\] sky130_fd_sc_hd__dfrtp_1
X_10996_ _05248_ _05251_ _05253_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ clknet_leaf_157_clk _00202_ net1140 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11622__S net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12666_ clknet_leaf_133_clk _00133_ net1196 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10746__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14405_ clknet_leaf_41_clk total_design.core.data_out_INSTR\[0\] net1092 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11617_ _05651_ net1746 net137 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10238__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09613__A1 total_design.core.data_cpu_o\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12597_ clknet_leaf_160_clk _00064_ net1142 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08216__B net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11420__A1 _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14336_ clknet_leaf_52_clk _01497_ net1094 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[27\]
+ sky130_fd_sc_hd__dfrtp_2
X_11548_ net1573 _05646_ net148 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06978__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold508 total_design.data_in_BUS\[15\] vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
X_14267_ clknet_leaf_46_clk _01446_ net1088 vssd1 vssd1 vccd1 vccd1 total_design.bus_full
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12453__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold519 total_design.lcd_display.row_1\[62\] vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
X_11479_ net1623 _05648_ net153 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13218_ clknet_leaf_126_clk _00685_ net1197 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14198_ clknet_leaf_112_clk _01378_ net1225 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_111_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ clknet_leaf_12_clk _00616_ net1025 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09762__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1208 total_design.core.regFile.register\[4\]\[10\] vssd1 vssd1 vccd1 vccd1 net2524
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 total_design.core.regFile.register\[21\]\[10\] vssd1 vssd1 vccd1 vccd1 net2535
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07710_ total_design.core.regFile.register\[22\]\[22\] net675 net578 total_design.core.regFile.register\[27\]\[22\]
+ _03218_ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08690_ _03958_ _03963_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__nor2_1
XANTENNA__10701__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ total_design.core.regFile.register\[14\]\[21\] net862 net807 total_design.core.regFile.register\[5\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__a22o_1
XANTENNA__06902__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07572_ _03044_ _03088_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09311_ _04194_ _04552_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__nor2_1
X_06523_ total_design.core.regFile.register\[9\]\[0\] net663 _02053_ _02090_ _02043_
+ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11532__S net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09242_ net318 _04261_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__nor2_1
XANTENNA__07863__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06454_ _01918_ _02020_ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_157_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09173_ _02439_ net447 net289 _04418_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10148__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06385_ net921 net948 net910 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout224_A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08124_ total_design.core.regFile.register\[9\]\[31\] net851 net835 total_design.core.regFile.register\[10\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__a22o_1
XANTENNA__09937__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06969__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ _03536_ _03537_ _03548_ _03549_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__or4_2
XFILLER_0_102_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1133_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07006_ total_design.core.regFile.register\[5\]\[9\] net630 net579 total_design.core.regFile.register\[27\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__a22o_1
XANTENNA__09368__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11487__B _05478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06214__X _01793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13756__Q total_design.core.data_bus_o\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout593_A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08040__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07394__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09525__X _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout760_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ _02187_ net508 net447 _02186_ _04209_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__o221a_1
XANTENNA__13193__RESET_B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_X net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11478__A1 _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10611__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ total_design.core.regFile.register\[21\]\[26\] net598 net567 total_design.core.regFile.register\[12\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__a22o_1
X_08888_ _04135_ _04141_ net324 vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__mux2_1
XANTENNA__07146__A2 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07839_ total_design.core.regFile.register\[20\]\[25\] net816 net815 total_design.core.regFile.register\[4\]\[25\]
+ net692 vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ _05096_ _05098_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_6_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09509_ _03184_ _04723_ _04741_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ total_design.core.data_bus_o\[21\] total_design.core.data_bus_o\[25\] total_design.core.data_bus_o\[29\]
+ net696 vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11442__S net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12520_ net976 net965 net882 _01714_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07854__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12451_ net2185 net206 net344 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10058__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11402_ _05593_ _05599_ _05472_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09847__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07606__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12382_ _01641_ _01642_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14121_ clknet_leaf_97_clk _01301_ net1246 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11333_ _05534_ _05529_ _05448_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_10_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14052_ clknet_leaf_100_clk _01232_ net1230 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11264_ _05432_ _05514_ _05520_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13003_ clknet_leaf_107_clk _00470_ net1224 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10215_ _04782_ net391 _04998_ vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08031__B1 _01992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11195_ _05449_ _05453_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__nand2_1
X_10146_ net185 net1933 net400 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__mux2_1
XANTENNA__11617__S net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11469__A1 _05655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10521__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10077_ net193 net2528 net406 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__mux2_1
XANTENNA__07137__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12130__A2 _05810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14497__Q total_design.core.ctrl.instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13905_ clknet_leaf_97_clk _01085_ net1245 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[115\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_195_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_195_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkload2_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13836_ clknet_leaf_59_clk _01044_ net1126 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10757__A _01771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13767_ clknet_leaf_58_clk total_design.core.data_mem.stored_data_adr\[10\] net1125
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[10\] sky130_fd_sc_hd__dfrtp_1
X_10979_ _05200_ _05202_ _05213_ _05199_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_139_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12448__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12718_ clknet_leaf_187_clk _00185_ net1031 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13698_ clknet_leaf_40_clk total_design.core.data_mem.stored_read_data\[5\] net1090
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_135_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12649_ clknet_leaf_17_clk _00116_ net1046 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09757__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06170_ total_design.core.data_cpu_o\[4\] vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold305 net80 vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14319_ clknet_leaf_67_clk _01480_ net1111 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold316 net89 vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 total_design.lcd_display.row_1\[100\] vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 total_design.lcd_display.row_2\[71\] vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold349 total_design.lcd_display.row_1\[73\] vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09860_ net254 net2762 net430 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__mux2_1
Xfanout807 net809 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_8
Xfanout818 _01968_ vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__clkbuf_8
Xfanout829 net830 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07376__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08811_ _02468_ net458 vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__and2_1
X_09791_ net254 total_design.core.regFile.register\[28\]\[10\] net438 vssd1 vssd1
+ vccd1 vccd1 _00113_ sky130_fd_sc_hd__mux2_1
Xhold1005 total_design.core.regFile.register\[26\]\[20\] vssd1 vssd1 vccd1 vccd1 net2321
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 total_design.core.regFile.register\[28\]\[27\] vssd1 vssd1 vccd1 vccd1 net2332
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ _03559_ _03602_ _03646_ _03997_ _02025_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__a41o_1
Xhold1027 total_design.core.regFile.register\[21\]\[16\] vssd1 vssd1 vccd1 vccd1 net2343
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10431__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1038 total_design.core.regFile.register\[18\]\[14\] vssd1 vssd1 vccd1 vccd1 net2354
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 total_design.core.regFile.register\[2\]\[4\] vssd1 vssd1 vccd1 vccd1 net2365
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07128__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12121__A2 _05804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09522__B1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08673_ total_design.keypad0.counter\[0\] total_design.keypad0.counter\[1\] total_design.keypad0.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_186_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_186_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07624_ _03136_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07555_ total_design.core.regFile.register\[10\]\[19\] net835 net765 total_design.core.regFile.register\[6\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__a22o_1
XANTENNA__08089__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout341_A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1083_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout439_A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06506_ net740 net739 net723 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__and3_1
XANTENNA__07836__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07486_ total_design.core.regFile.register\[11\]\[18\] net612 net608 total_design.core.regFile.register\[18\]\[18\]
+ _03006_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__a221o_1
XANTENNA__07300__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09225_ total_design.core.math.pc_val\[8\] _04448_ vssd1 vssd1 vccd1 vccd1 _04471_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06583__C net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06437_ total_design.core.ctrl.instruction\[0\] total_design.core.ctrl.instruction\[1\]
+ total_design.core.ctrl.instruction\[2\] vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout606_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout227_X net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09156_ _02390_ _02441_ _04403_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06368_ total_design.core.regFile.register\[14\]\[0\] net922 net917 net947 vssd1
+ vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__and4_1
XANTENNA__10199__A1 _04474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08107_ _03598_ _03599_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__nand2_2
XANTENNA__10606__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09087_ net463 _04229_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__nor2_1
X_06299_ total_design.core.instr_mem.instruction_adr_i\[1\] total_design.core.instr_mem.instruction_adr_stored\[1\]
+ net984 vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_110_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08038_ total_design.core.regFile.register\[13\]\[29\] net666 net562 total_design.core.regFile.register\[3\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold850 total_design.core.regFile.register\[23\]\[2\] vssd1 vssd1 vccd1 vccd1 net2166
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 total_design.core.regFile.register\[25\]\[10\] vssd1 vssd1 vccd1 vccd1 net2177
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold872 total_design.core.regFile.register\[6\]\[15\] vssd1 vssd1 vccd1 vccd1 net2188
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 total_design.core.regFile.register\[11\]\[28\] vssd1 vssd1 vccd1 vccd1 net2199
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 total_design.core.regFile.register\[25\]\[17\] vssd1 vssd1 vccd1 vccd1 net2210
+ sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ net234 net2006 net415 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__mux2_1
XANTENNA__13863__D total_design.core.ctrl.imm_32\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ net268 net2826 net414 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__S net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10341__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07119__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1550 net86 vssd1 vssd1 vccd1 vccd1 net2866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1561 total_design.core.regFile.register\[12\]\[1\] vssd1 vssd1 vccd1 vccd1 net2877
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout930_X net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ _05732_ _05742_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_177_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_177_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11961__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10902_ _05139_ _05145_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_28_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06477__D net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11882_ net897 _02118_ _05761_ _05762_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_28_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10833_ _05076_ _05082_ _05091_ _05080_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__a2bb2o_1
X_13621_ clknet_leaf_52_clk net1319 net1100 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06774__B total_design.core.ctrl.imm_32\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10764_ _01870_ _05022_ _01859_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__mux2_1
X_13552_ clknet_leaf_182_clk _01019_ net1040 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07827__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09292__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12503_ net974 total_design.core.instr_mem.instruction_i\[15\] vssd1 vssd1 vccd1
+ vccd1 _01706_ sky130_fd_sc_hd__and2b_1
X_13483_ clknet_leaf_108_clk _00950_ net1204 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10695_ net269 net2093 net358 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__mux2_1
X_12434_ net2539 net271 net345 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12365_ _01615_ _01624_ _01625_ _01627_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_101_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10516__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11201__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11316_ _05566_ _05567_ _05574_ net294 vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__a211oi_1
X_14104_ clknet_leaf_99_clk _01284_ net1229 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_12296_ _06131_ _06132_ _06133_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14035_ clknet_leaf_89_clk _01215_ net1260 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08213__C _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11247_ _05498_ _05504_ _05408_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08004__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ _05434_ _05436_ _05431_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10251__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10129_ net263 total_design.core.regFile.register\[18\]\[8\] net401 vssd1 vssd1 vccd1
+ vccd1 _00431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12103__A2 _05826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_168_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_168_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_106_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07530__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13819_ clknet_leaf_71_clk total_design.core.data_mem.data_cpu_i\[28\] net1206 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07340_ total_design.core.regFile.register\[15\]\[15\] net848 net766 total_design.core.regFile.register\[6\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07271_ total_design.core.regFile.register\[4\]\[14\] net623 net580 total_design.core.regFile.register\[27\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09010_ net335 _03596_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__nor2_1
X_06222_ total_design.core.instr_mem.instruction_adr_i\[14\] total_design.core.instr_mem.instruction_adr_stored\[14\]
+ net983 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__mux2_1
XANTENNA__09487__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06153_ total_design.core.ctrl.instruction\[20\] vssd1 vssd1 vccd1 vccd1 _01736_
+ sky130_fd_sc_hd__inv_2
XANTENNA__10426__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold102 total_design.core.instr_mem.instruction_adr_stored\[9\] vssd1 vssd1 vccd1
+ vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold113 total_design.core.data_mem.data_bus_i_reg\[1\] vssd1 vssd1 vccd1 vccd1 net1429
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 total_design.core.data_mem.data_read_adr_reg2\[26\] vssd1 vssd1 vccd1 vccd1
+ net1440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 total_design.core.instr_mem.instruction_adr_stored\[10\] vssd1 vssd1 vccd1
+ vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold146 total_design.core.data_mem.data_read_adr_reg2\[29\] vssd1 vssd1 vccd1 vccd1
+ net1462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold157 total_design.core.data_mem.data_cpu_i_reg\[5\] vssd1 vssd1 vccd1 vccd1 net1473
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 total_design.core.data_mem.data_cpu_i_reg\[24\] vssd1 vssd1 vccd1 vccd1 net1484
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09912_ net173 net2313 net428 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__mux2_1
Xhold179 total_design.core.data_mem.data_bus_i_reg\[30\] vssd1 vssd1 vccd1 vccd1 net1495
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout604 net607 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_8
Xfanout615 _02070_ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_4
XANTENNA__07349__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout626 net627 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_4
Xfanout637 net638 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__buf_4
X_09843_ net176 net2430 net436 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__mux2_1
Xfanout648 net649 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__clkbuf_8
Xfanout659 net662 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout389_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10161__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06986_ _02535_ _02515_ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__nand2b_1
X_09774_ net184 total_design.core.regFile.register\[29\]\[26\] net444 vssd1 vssd1
+ vccd1 vccd1 _00097_ sky130_fd_sc_hd__mux2_1
X_08725_ _03982_ _03983_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_159_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_159_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_174_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08656_ _03939_ net712 _03938_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__and3b_1
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07607_ total_design.core.regFile.register\[26\]\[20\] net869 net831 total_design.core.regFile.register\[31\]\[20\]
+ _03117_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09251__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _03860_ net880 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[8\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout344_X net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07538_ total_design.core.regFile.register\[23\]\[19\] net679 _03053_ _03055_ net687
+ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__a2111o_1
XANTENNA_clkbuf_leaf_189_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07469_ _02990_ _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__nand2_2
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout609_X net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09208_ _02491_ _04428_ _04453_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__a21o_1
X_10480_ net209 net2510 net378 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07037__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ _04384_ _04387_ net319 vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12030__A1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10336__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07588__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ total_design.lcd_display.row_2\[95\] _05837_ _05845_ total_design.lcd_display.row_2\[23\]
+ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11101_ net516 _05062_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__nand2_2
X_12081_ total_design.lcd_display.row_2\[108\] _05834_ _05852_ total_design.lcd_display.row_2\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__a22o_1
Xhold680 total_design.core.regFile.register\[24\]\[7\] vssd1 vssd1 vccd1 vccd1 net1996
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_127_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold691 total_design.core.regFile.register\[4\]\[25\] vssd1 vssd1 vccd1 vccd1 net2007
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ total_design.core.data_bus_o\[0\] net696 vssd1 vssd1 vccd1 vccd1 _05291_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_34_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10071__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07760__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06488__C net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ clknet_leaf_123_clk _00450_ net1186 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08984__B _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1380 total_design.core.regFile.register\[21\]\[24\] vssd1 vssd1 vccd1 vccd1 net2696
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1391 total_design.core.regFile.register\[30\]\[11\] vssd1 vssd1 vccd1 vccd1 net2707
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11934_ total_design.keypad0.key_out\[14\] net529 net475 total_design.keypad0.key_out\[10\]
+ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06785__A total_design.core.ctrl.instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07512__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11865_ total_design.lcd_display.currentState\[5\] _05748_ vssd1 vssd1 vccd1 vccd1
+ _05749_ sky130_fd_sc_hd__and2b_2
XFILLER_0_19_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13604_ clknet_leaf_62_clk net1336 net1125 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10816_ _05058_ _05061_ _05068_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__or3b_1
XFILLER_0_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11796_ net713 net1686 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_60_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13535_ clknet_leaf_156_clk _01002_ net1140 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_153_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10747_ total_design.core.regFile.register\[0\]\[22\] net355 vssd1 vssd1 vccd1 vccd1
+ _01021_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11630__S net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10280__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10678_ net211 net2351 net362 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13466_ clknet_leaf_124_clk _00933_ net1186 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09017__A2 _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10754__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12417_ _01672_ _01673_ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10246__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13397_ clknet_leaf_157_clk _00864_ net1141 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13225__RESET_B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12348_ _01612_ total_design.core.math.pc_val\[22\] net522 vssd1 vssd1 vccd1 vccd1
+ _01492_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06251__A2 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10770__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ net993 _04633_ net895 vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12461__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09725__B1 _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ clknet_leaf_87_clk _01198_ net1248 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06840_ total_design.core.ctrl.instruction\[26\] _02345_ vssd1 vssd1 vccd1 vccd1
+ _02398_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_108_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07200__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09770__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07751__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12860__RESET_B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06771_ _02318_ _02319_ _02331_ _02332_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__or4_1
X_08510_ total_design.keypad0.key_out\[10\] total_design.keypad0.key_out\[8\] _03717_
+ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09490_ _03136_ _04722_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_19_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07503__A2 _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ _03767_ _03795_ _03770_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_19_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06711__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08372_ _03725_ _03729_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_173_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11599__A0 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_944 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07323_ total_design.core.regFile.register\[21\]\[15\] net599 net564 total_design.core.regFile.register\[3\]\[15\]
+ _02850_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11540__S net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout137_A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07254_ net552 total_design.core.data_mem.data_cpu_i\[13\] total_design.core.ctrl.imm_32\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06205_ total_design.core.data_adr_o\[18\] _01783_ net962 vssd1 vssd1 vccd1 vccd1
+ _01784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10156__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07185_ total_design.core.regFile.register\[10\]\[12\] net837 net782 total_design.core.regFile.register\[27\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1046_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09945__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout401 _04990_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_4
XANTENNA__07990__A2 _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout412 net413 vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07318__X total_design.core.ctrl.imm_32\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout423 net425 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_6
Xfanout434 _04973_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout445 _04969_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__buf_4
Xfanout456 _04117_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_4
X_09826_ net255 net2032 net434 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__mux2_1
Xfanout467 net468 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_2
Xfanout478 net479 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_8
Xfanout489 net490 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_6
XANTENNA__07742__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ net251 net2656 net445 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__mux2_1
X_06969_ total_design.core.regFile.register\[8\]\[8\] net804 _02516_ _02519_ vssd1
+ vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout938_A _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout559_X net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06950__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ total_design.keypad0.counter\[3\] total_design.keypad0.counter\[5\] total_design.keypad0.counter\[7\]
+ total_design.keypad0.counter\[2\] vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__or4bb_1
X_09688_ _03557_ _04911_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__nand2_1
XANTENNA__09495__A2 _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08639_ _03924_ _03926_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_81_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11650_ _05651_ net1647 net133 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10601_ net262 net2630 net367 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__mux2_1
X_11581_ _05646_ net1694 net143 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09652__C1 _04100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11450__S net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10532_ net260 net2168 net376 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__mux2_1
X_13320_ clknet_leaf_171_clk _00787_ net1056 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10463_ net276 net1937 net377 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__mux2_1
X_13251_ clknet_leaf_8_clk _00718_ net1018 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10066__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12202_ total_design.core.math.pc_val\[6\] net528 _06050_ vssd1 vssd1 vccd1 vccd1
+ _01476_ sky130_fd_sc_hd__a21o_1
XANTENNA__09855__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11957__Y _05819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13182_ clknet_leaf_175_clk _00649_ net1053 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10394_ _04974_ net532 vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__nand2_1
X_12133_ total_design.lcd_display.row_2\[110\] _05834_ _05977_ _05980_ _05988_ vssd1
+ vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_36_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07981__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ total_design.lcd_display.row_1\[3\] _05830_ _05853_ total_design.lcd_display.row_2\[115\]
+ _05913_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__a221o_1
X_14527__1299 vssd1 vssd1 vccd1 vccd1 net1299 _14527__1299/LO sky130_fd_sc_hd__conb_1
XANTENNA__06499__B net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ net520 _05271_ _05273_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_53_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07194__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout990 net992 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__buf_2
XANTENNA__07733__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11625__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12966_ clknet_leaf_200_clk _00433_ net1002 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10749__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _05793_ total_design.keypad0.key_out\[1\] net530 vssd1 vssd1 vccd1 vccd1
+ _01448_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ clknet_leaf_123_clk _00364_ net1167 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11848_ total_design.lcd_display.currentState\[0\] total_design.lcd_display.currentState\[2\]
+ _05722_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_173_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13477__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12456__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11779_ net1827 net954 _05699_ _01782_ vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13518_ clknet_leaf_190_clk _00985_ net1032 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14498_ clknet_leaf_33_clk _01565_ net1070 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[26\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkload11 clknet_leaf_196_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__inv_6
XFILLER_0_125_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13449_ clknet_leaf_16_clk _00916_ net1024 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload22 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__bufinv_16
Xclkload33 clknet_leaf_187_clk vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__clkinv_4
Xclkload44 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__inv_8
XFILLER_0_24_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09765__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload55 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_77_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload66 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload77 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_77_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09410__A2 _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload88 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__07957__C1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload99 clknet_leaf_153_clk vssd1 vssd1 vccd1 vccd1 clkload99/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__08889__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10704__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08990_ _04239_ _04242_ net463 vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__mux2_1
XANTENNA__07972__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07941_ total_design.core.data_mem.data_cpu_i\[27\] vssd1 vssd1 vccd1 vccd1 _03440_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_166_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09174__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07872_ _03373_ _03374_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__xor2_4
XANTENNA__07185__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ _04838_ _04839_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06823_ total_design.core.regFile.register\[18\]\[5\] net858 net835 total_design.core.regFile.register\[10\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06696__Y _02263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09542_ _03230_ net509 _04418_ _04664_ _04766_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__o221a_1
X_06754_ total_design.core.regFile.register\[22\]\[4\] net674 net624 total_design.core.regFile.register\[14\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07314__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06685_ total_design.core.regFile.register\[9\]\[3\] net851 net780 total_design.core.regFile.register\[27\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a22o_1
X_09473_ _04253_ _04257_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_90_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08424_ _03777_ _03778_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08355_ total_design.keypad0.key_out\[5\] total_design.keypad0.key_out\[7\] vssd1
+ vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__nand2_1
Xclkbuf_4_9__f_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1163_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07306_ net552 total_design.core.data_mem.data_cpu_i\[14\] total_design.core.ctrl.imm_32\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__a21oi_1
Xclkload5 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_73_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08286_ net1460 net941 _03677_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[0\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06999__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11992__B1 _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07237_ total_design.core.regFile.register\[20\]\[13\] net818 net790 total_design.core.regFile.register\[24\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07168_ total_design.core.regFile.register\[22\]\[12\] net677 net608 total_design.core.regFile.register\[18\]\[12\]
+ _02702_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout790_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10614__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07099_ total_design.core.ctrl.instruction\[30\] _02541_ total_design.core.ctrl.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08151__Y _03642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1207 net1210 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1218 net1219 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__clkbuf_4
Xfanout220 net223 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__clkbuf_2
Xfanout1229 net1231 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__clkbuf_4
Xfanout231 _04589_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
Xfanout253 net256 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_2
Xfanout264 _04475_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07176__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 _04426_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07715__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout286 net287 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_2
XANTENNA__09704__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09809_ net174 net2125 net439 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__mux2_1
Xfanout297 _04192_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout843_X net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06923__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11445__S net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ clknet_leaf_142_clk _00287_ net1176 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12751_ clknet_leaf_161_clk _00218_ net1151 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08140__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06485__D net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11702_ net6 net935 net878 net1796 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__o22a_1
X_12682_ clknet_leaf_20_clk _00149_ net1050 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14421_ clknet_leaf_29_clk total_design.core.data_out_INSTR\[16\] net1073 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[16\] sky130_fd_sc_hd__dfrtp_1
X_11633_ _05679_ net1704 net135 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14352_ clknet_leaf_45_clk _00021_ net1086 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06274__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11564_ _05667_ net1820 net141 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13303_ clknet_leaf_162_clk _00770_ net1166 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_98_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10515_ net203 net2350 net482 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11495_ net1570 _05627_ net151 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__mux2_1
X_14283_ net987 _01459_ net1083 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07894__A _03395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13234_ clknet_leaf_145_clk _00701_ net1179 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10446_ net218 net2271 net384 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13165_ clknet_leaf_0_clk _00632_ net1005 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10524__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10377_ net226 net2750 net487 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07954__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12116_ total_design.lcd_display.row_1\[38\] _05827_ _05838_ total_design.lcd_display.row_1\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__a22o_1
X_13096_ clknet_leaf_169_clk _00563_ net1159 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12047_ total_design.lcd_display.row_1\[2\] _05830_ _05904_ _05906_ vssd1 vssd1 vccd1
+ vccd1 _05907_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_144_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07167__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07706__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09614__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13998_ clknet_leaf_97_clk _01178_ net1246 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12949_ clknet_leaf_157_clk _00416_ net1140 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06395__D net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06470_ _01924_ net901 _02018_ _01742_ total_design.core.ctrl.instruction\[15\] vssd1
+ vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__o311a_1
XFILLER_0_157_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06693__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08140_ total_design.core.regFile.register\[14\]\[31\] net625 net583 total_design.core.regFile.register\[6\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload100 clknet_leaf_154_clk vssd1 vssd1 vccd1 vccd1 clkload100/Y sky130_fd_sc_hd__inv_8
X_08071_ total_design.core.regFile.register\[30\]\[30\] net840 net812 total_design.core.regFile.register\[23\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__a22o_1
Xclkload111 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 clkload111/Y sky130_fd_sc_hd__inv_6
Xclkload122 clknet_leaf_137_clk vssd1 vssd1 vccd1 vccd1 clkload122/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_116_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload133 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 clkload133/X sky130_fd_sc_hd__clkbuf_4
X_07022_ total_design.core.regFile.register\[20\]\[9\] net817 net766 total_design.core.regFile.register\[6\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a22o_1
XANTENNA__12518__A2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload144 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 clkload144/X sky130_fd_sc_hd__clkbuf_8
Xclkload155 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 clkload155/Y sky130_fd_sc_hd__inv_6
XFILLER_0_114_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload166 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 clkload166/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_168_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload177 clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 clkload177/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_168_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09395__A1 total_design.core.ctrl.instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10434__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ net336 _02718_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__or2_1
Xhold17 total_design.core.data_mem.data_read_adr_reg\[26\] vssd1 vssd1 vccd1 vccd1
+ net1333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold28 total_design.core.data_mem.data_read_adr_reg\[0\] vssd1 vssd1 vccd1 vccd1
+ net1344 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ total_design.core.regFile.register\[18\]\[27\] net858 net851 total_design.core.regFile.register\[9\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__a22o_1
Xhold39 total_design.core.math.pc_val\[7\] vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12151__B1 _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1009_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ total_design.core.regFile.register\[23\]\[25\] net679 net583 total_design.core.regFile.register\[6\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout371_A _05013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06905__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06806_ _02359_ _02361_ _02363_ _02365_ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__or4_1
X_07786_ total_design.core.regFile.register\[9\]\[24\] net851 net811 total_design.core.regFile.register\[23\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__a22o_1
XANTENNA__06586__C net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07044__A total_design.core.ctrl.instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09525_ total_design.core.ctrl.instruction\[21\] net885 net754 total_design.core.data_cpu_o\[21\]
+ _04757_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__a221o_2
X_06737_ total_design.core.regFile.register\[30\]\[4\] net838 net783 total_design.core.regFile.register\[2\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_63_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout636_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08122__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06668_ net554 _02211_ _02235_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__a21o_1
X_09456_ _04691_ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08407_ net933 _03742_ _03741_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_136_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06684__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout803_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10609__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06599_ total_design.core.regFile.register\[29\]\[1\] net655 _02162_ _02165_ _02167_
+ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ _04625_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__inv_2
X_14526__1298 vssd1 vssd1 vccd1 vccd1 net1298 _14526__1298/LO sky130_fd_sc_hd__conb_1
XFILLER_0_164_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08338_ net1440 net938 _03703_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[26\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11013__B _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06436__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08269_ net1402 net557 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[19\]
+ sky130_fd_sc_hd__and2_1
X_10300_ net281 net2258 net492 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ _05481_ _05499_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10231_ net246 net1714 net500 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__mux2_1
XANTENNA__10344__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07397__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10162_ net265 net2743 net394 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout960_X net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1004 net1006 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__clkbuf_4
Xfanout1015 net1027 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1026 net1027 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_4
Xfanout1037 net1045 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10093_ net273 net2729 net404 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__mux2_1
Xfanout1048 net1051 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12142__B1 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 net1135 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13921_ clknet_leaf_97_clk _01101_ net1244 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09434__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06410__X _01986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13852_ clknet_leaf_52_clk _01060_ net1094 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09153__B _04401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06269__S net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11970__Y _05832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12803_ clknet_leaf_6_clk _00270_ net1017 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13783_ clknet_leaf_50_clk total_design.core.data_mem.stored_data_adr\[26\] net1100
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[26\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_54_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10995_ _05253_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__inv_2
XANTENNA__13069__RESET_B net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08113__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ clknet_leaf_174_clk _00201_ net1053 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07321__B1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06675__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12665_ clknet_leaf_197_clk _00132_ net1007 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10519__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08056__Y _03551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10208__A0 _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14404_ clknet_leaf_51_clk net1799 net1097 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11616_ _05650_ net1738 net139 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09613__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12596_ clknet_leaf_142_clk _00063_ net1175 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14335_ clknet_leaf_52_clk _01496_ net1094 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06427__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11547_ net1512 _05645_ net145 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold509 total_design.data_in_BUS\[7\] vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
X_14266_ clknet_leaf_63_clk _01445_ net1122 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_11478_ net1574 _05628_ net156 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13217_ clknet_leaf_121_clk _00684_ net1170 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10254__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10429_ net245 net2206 net381 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14197_ clknet_leaf_111_clk _01377_ net1225 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_2
XANTENNA__07388__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08232__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07927__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ clknet_leaf_28_clk _00615_ net1075 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ clknet_leaf_164_clk _00546_ net1164 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1209 total_design.core.regFile.register\[22\]\[19\] vssd1 vssd1 vccd1 vccd1 net2525
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08352__A2 _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07640_ total_design.core.regFile.register\[31\]\[21\] net832 net787 total_design.core.regFile.register\[13\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07560__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07571_ _03085_ _03086_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__nand2_2
XFILLER_0_48_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_45_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08104__A2 total_design.core.data_mem.data_cpu_i\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_06522_ total_design.core.regFile.register\[23\]\[0\] net681 _02041_ _02047_ _02095_
+ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__a2111o_1
X_09310_ _04366_ _04551_ net317 vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06453_ net973 _02025_ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__or2_1
X_09241_ _04194_ _04485_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10429__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09172_ net968 _02439_ _02440_ net537 vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_56_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06384_ total_design.core.regFile.register\[31\]\[0\] net927 net912 net947 vssd1
+ vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__nand4_1
XFILLER_0_56_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ total_design.core.regFile.register\[1\]\[31\] net828 _03611_ _03612_ _03614_
+ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout217_A _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08054_ total_design.core.regFile.register\[25\]\[29\] net647 net597 total_design.core.regFile.register\[21\]\[29\]
+ _03539_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14280__RESET_B net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07005_ total_design.core.regFile.register\[14\]\[9\] net626 _02552_ vssd1 vssd1
+ vccd1 vccd1 _02553_ sky130_fd_sc_hd__a21o_1
XANTENNA__10164__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11487__C _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07379__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07039__A _02564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09953__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout586_A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _02183_ net462 net504 vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__a21o_1
X_07907_ total_design.core.regFile.register\[2\]\[26\] net637 net634 total_design.core.regFile.register\[16\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ _04138_ _04140_ net459 vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__mux2_1
X_07838_ total_design.core.regFile.register\[16\]\[25\] net855 _03338_ _03339_ _03341_
+ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_169_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07551__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout920_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ _03275_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_36_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09508_ _03112_ _03133_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__nand2_1
X_10780_ total_design.core.data_bus_o\[16\] total_design.core.data_bus_o\[20\] total_design.core.data_bus_o\[23\]
+ total_design.core.data_bus_o\[31\] net696 vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__o41a_1
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09439_ total_design.core.math.pc_val\[17\] _04651_ vssd1 vssd1 vccd1 vccd1 _04676_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06657__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10339__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12450_ net2276 net210 net345 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11401_ _05651_ _05652_ _05655_ _05659_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__and4_1
XFILLER_0_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12381_ _01631_ _01632_ _01633_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08803__B1 total_design.core.data_mem.data_cpu_i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10610__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ clknet_leaf_111_clk _01300_ net1225 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11332_ _05530_ _05537_ _05448_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__a21o_1
XANTENNA__07082__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14051_ clknet_leaf_90_clk _01231_ net1261 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10074__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11263_ _05514_ _05520_ _05432_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_91_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07909__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13002_ clknet_leaf_19_clk _00469_ net1050 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11965__Y _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10214_ net1916 net392 vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__nand2_1
X_11194_ _05440_ _05442_ _05447_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__nand3_1
XFILLER_0_101_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08987__B _02367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10145_ net192 net2633 net400 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10076_ net197 net2462 net407 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__mux2_1
XANTENNA__08334__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13904_ clknet_leaf_74_clk _01084_ net1220 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07542__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13835_ clknet_leaf_58_clk _01043_ net1127 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06896__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11633__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13766_ clknet_leaf_58_clk total_design.core.data_mem.stored_data_adr\[9\] net1125
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09295__B1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10978_ _05236_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_139_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07412__A _02917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12717_ clknet_leaf_3_clk _00184_ net1014 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06648__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10249__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13697_ clknet_leaf_40_clk total_design.core.data_mem.stored_read_data\[4\] net1092
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12648_ clknet_leaf_170_clk _00115_ net1159 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_154_Left_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09598__A1 _03375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10773__A total_design.core.data_bus_o\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12579_ clknet_leaf_8_clk _00046_ net1017 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14318_ clknet_leaf_66_clk _01479_ net1122 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_123_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07073__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 total_design.lcd_display.row_1\[67\] vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold317 _01380_ vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold328 total_design.lcd_display.row_2\[91\] vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold339 total_design.lcd_display.row_2\[78\] vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06820__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14249_ clknet_leaf_109_clk _01429_ net1240 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09773__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout808 net809 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__buf_4
Xfanout819 net822 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08897__B _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08810_ net311 total_design.core.data_mem.data_cpu_i\[6\] vssd1 vssd1 vccd1 vccd1
+ _04065_ sky130_fd_sc_hd__nor2_1
XANTENNA__10712__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ net250 net2236 net440 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__mux2_1
XANTENNA__12106__B1 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1006 total_design.core.regFile.register\[30\]\[3\] vssd1 vssd1 vccd1 vccd1 net2322
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07781__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_163_Left_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1017 total_design.core.regFile.register\[19\]\[13\] vssd1 vssd1 vccd1 vccd1 net2333
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14525__1297 vssd1 vssd1 vccd1 vccd1 net1297 _14525__1297/LO sky130_fd_sc_hd__conb_1
X_08741_ _03375_ _03421_ _03512_ _03996_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__and4_1
Xhold1028 total_design.core.regFile.register\[13\]\[28\] vssd1 vssd1 vccd1 vccd1 net2344
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 total_design.core.regFile.register\[8\]\[17\] vssd1 vssd1 vccd1 vccd1 net2355
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08672_ net711 _03948_ _03949_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__and3_1
XANTENNA__07533__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07623_ _03134_ _03135_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__and2_2
XFILLER_0_89_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_18_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13895__CLK clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07554_ total_design.core.regFile.register\[23\]\[19\] net811 net799 total_design.core.regFile.register\[29\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06505_ total_design.core.regFile.register\[21\]\[0\] net747 net734 net729 vssd1
+ vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__and4_1
XFILLER_0_146_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07485_ total_design.core.regFile.register\[19\]\[18\] net640 net616 total_design.core.regFile.register\[10\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__a22o_1
XANTENNA__10159__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout334_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_172_Left_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09224_ _04457_ _04469_ _04124_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09948__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06436_ total_design.core.regFile.register\[0\]\[0\] net874 _02006_ _02011_ vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[0\] sky130_fd_sc_hd__o22a_4
XFILLER_0_63_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09155_ _02367_ _02389_ _04350_ _02341_ _04375_ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__a221o_1
X_06367_ net921 net916 net947 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout501_A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1243_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10199__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08106_ _03595_ _03597_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__or2_2
XANTENNA__07064__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06298_ total_design.core.data_mem.data_read net997 total_design.core.data_adr_o\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09086_ _04335_ _04336_ net328 vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__mux2_1
XANTENNA__08153__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08037_ _03532_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[29\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06811__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold840 total_design.core.regFile.register\[3\]\[5\] vssd1 vssd1 vccd1 vccd1 net2156
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11148__B2 _05358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold851 total_design.core.regFile.register\[22\]\[29\] vssd1 vssd1 vccd1 vccd1 net2167
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 total_design.core.regFile.register\[22\]\[11\] vssd1 vssd1 vccd1 vccd1 net2178
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 total_design.core.regFile.register\[6\]\[12\] vssd1 vssd1 vccd1 vccd1 net2189
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 total_design.core.regFile.register\[29\]\[17\] vssd1 vssd1 vccd1 vccd1 net2200
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 total_design.core.regFile.register\[4\]\[22\] vssd1 vssd1 vccd1 vccd1 net2211
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_X net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10622__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ net276 net2342 net414 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__mux2_1
X_08939_ _02338_ _04104_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08316__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09513__A1 _03187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1540 total_design.core.regFile.register\[5\]\[4\] vssd1 vssd1 vccd1 vccd1 net2856
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10659__A0 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1551 total_design.core.regFile.register\[12\]\[24\] vssd1 vssd1 vccd1 vccd1 net2867
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11950_ _05809_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__nor2_4
Xhold1562 total_design.core.regFile.register\[23\]\[17\] vssd1 vssd1 vccd1 vccd1 net2878
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10901_ _05157_ _05159_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09712__A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06878__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ total_design.core.math.pc_val\[0\] total_design.core.program_count.imm_val_reg\[0\]
+ _05760_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_28_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout923_X net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11453__S net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13620_ clknet_leaf_50_clk net1347 net1097 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10832_ _05076_ _05085_ _05079_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_45_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13551_ clknet_leaf_161_clk _01018_ net1151 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10763_ _01861_ _01869_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10069__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09858__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12502_ net974 total_design.core.ctrl.instruction\[14\] net881 _01705_ vssd1 vssd1
+ vccd1 vccd1 _01553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13482_ clknet_leaf_19_clk _00949_ net1049 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10694_ net278 net2533 net359 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12433_ net1900 net277 net345 vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__mux2_1
XANTENNA__07055__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12364_ net991 _01626_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_130_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14103_ clknet_leaf_98_clk _01283_ net1242 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_11315_ _05564_ _05565_ _05567_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06802__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12295_ total_design.core.math.pc_val\[17\] total_design.core.program_count.imm_val_reg\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09593__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14034_ clknet_leaf_88_clk _01214_ net1250 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[116\]
+ sky130_fd_sc_hd__dfrtp_1
X_11246_ _05498_ _05504_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11628__S net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10532__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ _05422_ _05423_ _05429_ _05433_ _05357_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__a311o_1
XFILLER_0_101_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07763__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10128_ net265 net2851 net398 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__mux2_1
XANTENNA__06311__A _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08307__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10059_ net258 net2716 net408 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__mux2_1
XANTENNA__07515__B1 total_design.core.ctrl.imm_32\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09622__A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12459__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06869__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13818_ clknet_leaf_71_clk total_design.core.data_mem.data_cpu_i\[27\] net1206 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13749_ clknet_leaf_73_clk total_design.core.data_mem.stored_write_data\[24\] net1209
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[24\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_174_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09768__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07270_ total_design.core.regFile.register\[20\]\[14\] net673 net581 total_design.core.regFile.register\[6\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__a22o_1
XANTENNA__07294__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06221_ total_design.core.data_adr_o\[8\] _01799_ net963 vssd1 vssd1 vccd1 vccd1
+ _01800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10707__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06152_ total_design.core.ctrl.instruction\[3\] vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__inv_2
Xhold103 total_design.core.instr_mem.instruction_adr_stored\[22\] vssd1 vssd1 vccd1
+ vccd1 net1419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold114 total_design.core.instr_mem.instruction_adr_stored\[1\] vssd1 vssd1 vccd1
+ vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10790__X _05049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold125 total_design.core.instr_mem.instruction_adr_stored\[26\] vssd1 vssd1 vccd1
+ vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold136 total_design.core.math.pc_val\[22\] vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold147 total_design.core.data_mem.data_read_adr_reg2\[16\] vssd1 vssd1 vccd1 vccd1
+ net1463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold158 total_design.core.data_mem.data_bus_i_reg\[24\] vssd1 vssd1 vccd1 vccd1 net1474
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ net179 net2243 net428 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__mux2_1
Xhold169 total_design.core.math.pc_val\[17\] vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout605 net607 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11538__S net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout616 net619 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09743__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09842_ net183 net1958 net436 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__mux2_1
Xfanout627 _02064_ vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__buf_4
XANTENNA__10442__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout638 net639 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__buf_4
Xfanout649 net650 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11550__A1 _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07754__B1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ net188 net1980 net444 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__mux2_1
X_06985_ net555 total_design.core.data_mem.data_cpu_i\[8\] total_design.core.ctrl.imm_32\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout284_A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08724_ _01734_ net36 net38 net37 vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__or4_2
XANTENNA__07506__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08655_ total_design.lcd_display.cnt_500hz\[7\] total_design.lcd_display.cnt_500hz\[8\]
+ _03936_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout549_A total_design.core.data_mem.next_write vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_117_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07606_ total_design.core.regFile.register\[5\]\[20\] net806 net798 total_design.core.regFile.register\[29\]\[20\]
+ _03114_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__a221o_1
XANTENNA__09251__B _04495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08586_ _03842_ net880 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[7\]
+ sky130_fd_sc_hd__nor2_1
X_07537_ total_design.core.regFile.register\[26\]\[19\] net645 net609 total_design.core.regFile.register\[18\]\[19\]
+ _03054_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout337_X net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07285__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07468_ _02969_ _02989_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__or2_2
XFILLER_0_174_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ _02108_ net458 _02468_ _02448_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06419_ total_design.core.ctrl.instruction\[22\] total_design.core.ctrl.instruction\[24\]
+ net918 _01936_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__and4_4
XFILLER_0_107_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout504_X net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10617__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__A1 total_design.core.data_bus_o\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07399_ total_design.core.regFile.register\[30\]\[16\] net839 net817 total_design.core.regFile.register\[20\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__a22o_1
XANTENNA__07037__A2 total_design.core.data_mem.data_cpu_i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09138_ _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__inv_2
XANTENNA__12030__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06340__A_N total_design.core.ctrl.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__06245__A0 total_design.core.instr_mem.instruction_adr_i\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09069_ _02292_ net705 _04319_ net536 vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11100_ net516 _05078_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__nand2_2
XFILLER_0_130_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07993__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ total_design.lcd_display.row_1\[68\] _05804_ _05848_ total_design.lcd_display.row_2\[124\]
+ _05937_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 total_design.core.regFile.register\[22\]\[0\] vssd1 vssd1 vccd1 vccd1 net1986
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 total_design.core.regFile.register\[7\]\[3\] vssd1 vssd1 vccd1 vccd1 net1997
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11448__S net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold692 total_design.core.regFile.register\[20\]\[3\] vssd1 vssd1 vccd1 vccd1 net2008
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ _05287_ _05288_ _05289_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a21o_1
XANTENNA__10352__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__A1 _05636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12097__A2 _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ clknet_leaf_156_clk _00449_ net1140 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1370 total_design.core.regFile.register\[18\]\[1\] vssd1 vssd1 vccd1 vccd1 net2686
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1381 total_design.core.regFile.register\[4\]\[18\] vssd1 vssd1 vccd1 vccd1 net2697
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07514__X total_design.core.data_mem.data_cpu_i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ total_design.keypad0.key_out\[13\] net529 net475 net933 vssd1 vssd1 vccd1
+ vccd1 _01460_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1392 total_design.core.regFile.register\[22\]\[31\] vssd1 vssd1 vccd1 vccd1 net2708
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06277__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11864_ _01723_ _05722_ _05747_ total_design.lcd_display.currentState\[3\] vssd1
+ vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__a22o_1
XANTENNA__08058__A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13603_ clknet_leaf_60_clk net1340 net1132 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10815_ _05058_ _05061_ _05068_ _05073_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_89_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11795_ net1826 _01911_ _05694_ _01822_ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13534_ clknet_leaf_174_clk _01001_ net1054 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_10746_ net2014 net355 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07276__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09670__B1 _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14524__1296 vssd1 vssd1 vccd1 vccd1 net1296 _14524__1296/LO sky130_fd_sc_hd__conb_1
XFILLER_0_152_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13465_ clknet_leaf_197_clk _00932_ net1007 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10527__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10677_ net217 net2238 net361 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__mux2_1
XANTENNA__08064__Y _03559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12416_ total_design.core.math.pc_val\[30\] net989 vssd1 vssd1 vccd1 vccd1 _01673_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07028__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12021__A2 _05826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06306__A _01852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13396_ clknet_leaf_140_clk _00863_ net1183 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06236__A0 total_design.core.instr_mem.instruction_adr_i\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12347_ net899 _03234_ _01611_ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06833__A_N _02367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07984__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12278_ _06114_ _06116_ _06113_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10770__B _05028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14017_ clknet_leaf_96_clk _01197_ net1253 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09725__A1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ _05484_ _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11532__A1 _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08240__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07736__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07200__A2 total_design.core.data_mem.data_cpu_i\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12088__A2 _05814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ total_design.core.regFile.register\[9\]\[4\] net663 net566 total_design.core.regFile.register\[12\]\[4\]
+ _02321_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__a221o_1
XANTENNA__10769__Y _05028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08440_ _03792_ _03793_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_19_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire305_X net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08371_ total_design.keypad0.key_out\[8\] _03728_ vssd1 vssd1 vccd1 vccd1 _03729_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07322_ total_design.core.regFile.register\[13\]\[15\] net668 net638 total_design.core.regFile.register\[2\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07267__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09661__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07253_ _02776_ _02782_ _02788_ _02771_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[13\]
+ sky130_fd_sc_hd__o31a_4
XFILLER_0_45_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10437__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06204_ total_design.core.instr_mem.instruction_adr_i\[18\] total_design.core.instr_mem.instruction_adr_stored\[18\]
+ net981 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07184_ total_design.core.regFile.register\[9\]\[12\] net852 net818 total_design.core.regFile.register\[20\]\[12\]
+ _02722_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a221o_1
XANTENNA__07019__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12012__A2 _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10961__A total_design.core.data_bus_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1039_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09527__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout499_A _05004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 net405 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_6
XANTENNA__10172__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout413 _04985_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_4
XANTENNA__09716__B2 _04604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09246__B _04102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout424 net425 vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1206_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11523__A1 _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07727__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 _04973_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09961__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout446 _04189_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ net249 net2684 net437 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__mux2_1
Xfanout468 _02184_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_2
XANTENNA_fanout666_A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 _05015_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_4
XANTENNA_fanout287_X net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ net261 net2849 net445 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__mux2_1
XANTENNA__12079__A2 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06968_ total_design.core.regFile.register\[2\]\[8\] net785 _02517_ _02518_ vssd1
+ vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__a211o_1
X_08707_ total_design.keypad0.counter\[4\] _03951_ vssd1 vssd1 vccd1 vccd1 _03972_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09687_ _04911_ _03557_ _04892_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__or3b_1
X_06899_ total_design.core.regFile.register\[11\]\[7\] net615 net566 total_design.core.regFile.register\[12\]\[7\]
+ _02452_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout833_A _01959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08152__B1 total_design.core.ctrl.imm_32\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08638_ _03924_ _03926_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__and2_1
XANTENNA_hold244_A total_design.core.math.pc_val\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06702__A1 _02213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07988__Y _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_0__f_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout621_X net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ net2882 net340 net718 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[24\]
+ sky130_fd_sc_hd__and3_1
X_10600_ net266 net2411 net365 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__mux2_1
X_11580_ _05645_ net1828 net141 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13869__D total_design.core.ctrl.imm_32\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10531_ net282 net2379 net373 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10347__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07663__C1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13250_ clknet_leaf_130_clk _00717_ net1199 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12003__A2 _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10462_ net244 net1884 net380 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__mux2_1
XANTENNA__09404__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12201_ net902 _02442_ _06049_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__a21oi_1
X_13181_ clknet_leaf_10_clk _00648_ net1019 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10393_ net161 net2858 net486 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__mux2_1
X_12132_ _05982_ _05984_ _05985_ _05987_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__or4_1
XANTENNA__11686__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07430__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12063_ total_design.lcd_display.row_2\[83\] _05818_ _05821_ total_design.lcd_display.row_1\[43\]
+ _05921_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__a221o_1
XANTENNA__10082__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11514__A1 _05645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09871__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ _05253_ _05256_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11973__Y _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06499__C net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09724__X _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08995__B _03322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout980 net985 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_2
Xfanout991 net992 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__buf_2
XANTENNA__09443__Y _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ clknet_leaf_113_clk _00432_ net1203 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08143__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11916_ _03908_ _05777_ _05786_ _01734_ _05792_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07497__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12490__A2 total_design.core.ctrl.instruction\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12896_ clknet_leaf_191_clk _00363_ net1032 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11847_ total_design.lcd_display.currentState\[0\] net709 _05733_ vssd1 vssd1 vccd1
+ vccd1 _01438_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14566_ net38 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07249__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11778_ net1836 net954 _05699_ _01802_ vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13517_ clknet_leaf_6_clk _00984_ net1017 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10729_ total_design.core.regFile.register\[0\]\[4\] net353 vssd1 vssd1 vccd1 vccd1
+ _01003_ sky130_fd_sc_hd__and2_1
XANTENNA__10257__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14497_ clknet_leaf_36_clk _01564_ net1070 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_70_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08235__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload12 clknet_leaf_197_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinv_4
X_13448_ clknet_leaf_24_clk _00915_ net1057 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload23 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__inv_6
XFILLER_0_140_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload34 clknet_leaf_188_clk vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_51_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_173_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload45 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload56 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__inv_12
Xclkload67 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__inv_12
X_13379_ clknet_leaf_5_clk _00846_ net1024 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload78 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_77_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11753__B2 total_design.core.data_bus_o\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload89 clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_149_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09159__C1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07940_ _03426_ _03427_ _03439_ net875 total_design.core.regFile.register\[0\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[27\] sky130_fd_sc_hd__o32a_4
XANTENNA_clkbuf_4_11__f_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_188_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09781__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09174__A2 _04410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07871_ _03323_ _03327_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__nand2_2
X_09610_ total_design.core.math.pc_val\[24\] _04799_ total_design.core.math.pc_val\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ total_design.core.regFile.register\[30\]\[5\] net840 net812 total_design.core.regFile.register\[23\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a22o_1
XANTENNA__10720__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ _04194_ _04771_ _04772_ _04410_ net295 vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__o32a_1
X_06753_ _02267_ _02290_ _02289_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08134__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07314__B _02845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09472_ net319 _04332_ _04666_ _04706_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a31o_1
XANTENNA__07488__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06684_ total_design.core.regFile.register\[31\]\[3\] net832 net791 total_design.core.regFile.register\[24\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08423_ _03773_ _03776_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11551__S net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_126_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08354_ total_design.keypad0.key_out\[13\] net931 total_design.keypad0.key_out\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07305_ _02821_ _02824_ _02837_ net874 total_design.core.regFile.register\[0\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[14\] sky130_fd_sc_hd__o32a_4
XFILLER_0_46_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08285_ total_design.core.data_mem.data_write_adr_reg\[0\] net549 net541 total_design.core.data_mem.data_read_adr_reg\[0\]
+ net945 vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__a221o_1
Xclkload6 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__inv_8
XFILLER_0_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10167__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout414_A _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1156_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07236_ total_design.core.regFile.register\[30\]\[13\] net838 net798 total_design.core.regFile.register\[29\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__a22o_1
XANTENNA__07660__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07167_ total_design.core.regFile.register\[25\]\[12\] net649 net625 total_design.core.regFile.register\[14\]\[12\]
+ _02703_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a221o_1
XANTENNA__07948__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11744__B2 total_design.core.data_bus_o\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08161__A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07098_ total_design.core.ctrl.instruction\[20\] total_design.core.ctrl.instruction\[30\]
+ _02541_ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout783_A _01986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1208 net1210 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__buf_2
Xfanout210 _04721_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_1
Xfanout1219 net1222 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__clkbuf_2
Xfanout221 net223 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_2
Xfanout232 net235 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_2
XANTENNA__09544__X _04776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout243 _04543_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_2
Xfanout254 net256 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout571_X net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_2
Xfanout276 net279 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ net178 net2332 net439 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__mux2_1
Xfanout287 _04201_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10630__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09704__B _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout298 _04159_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_4
X_14523__1295 vssd1 vssd1 vccd1 vccd1 net1295 _14523__1295/LO sky130_fd_sc_hd__conb_1
X_09739_ _03645_ net509 _04624_ _04667_ _04959_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__o221a_1
XANTENNA__08125__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout836_X net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_clk_X clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12750_ clknet_leaf_189_clk _00217_ net1030 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07479__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11680__A0 _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11701_ net5 net935 net878 net1563 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__o22a_1
XFILLER_0_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12681_ clknet_leaf_16_clk _00148_ net1023 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11461__S net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14420_ clknet_leaf_31_clk total_design.core.data_out_INSTR\[15\] net1062 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[15\] sky130_fd_sc_hd__dfrtp_1
X_11632_ _05632_ net1791 net135 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14351_ clknet_leaf_45_clk _00038_ net1086 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11563_ _05665_ net1687 net141 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10077__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13302_ clknet_leaf_152_clk _00769_ net1139 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09866__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10514_ net206 net1985 net480 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__mux2_1
X_14282_ net987 _01458_ net1082 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11968__Y _05830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11494_ net1602 _05677_ net149 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__mux2_1
XANTENNA__07651__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13233_ clknet_leaf_152_clk _00700_ net1146 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10445_ _04681_ net2346 net381 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11735__B2 total_design.core.data_bus_o\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07403__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13164_ clknet_leaf_118_clk _00631_ net1169 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10376_ net235 net2744 net485 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12115_ _03928_ _05970_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__or2_1
X_13095_ clknet_leaf_174_clk _00562_ net1054 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12046_ total_design.lcd_display.row_2\[58\] _05835_ _05843_ total_design.lcd_display.row_1\[122\]
+ _05905_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_144_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11636__S net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10540__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09614__B _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13997_ clknet_leaf_91_clk _01177_ net1262 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12948_ clknet_leaf_141_clk _00415_ net1182 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11671__A0 _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06678__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10776__A total_design.core.data_bus_o\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12879_ clknet_leaf_161_clk _00346_ net1151 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07890__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07150__A _02666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10226__A1 _04966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14549_ net1269 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XANTENNA__09631__A3 _04296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09776__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08070_ total_design.core.regFile.register\[26\]\[30\] net871 net848 total_design.core.regFile.register\[15\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload101 clknet_leaf_155_clk vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_15_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07642__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload112 clknet_leaf_162_clk vssd1 vssd1 vccd1 vccd1 clkload112/Y sky130_fd_sc_hd__inv_6
XFILLER_0_71_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload123 clknet_leaf_138_clk vssd1 vssd1 vccd1 vccd1 clkload123/Y sky130_fd_sc_hd__inv_6
XFILLER_0_71_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload134 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 clkload134/Y sky130_fd_sc_hd__clkinvlp_4
X_07021_ total_design.core.regFile.register\[25\]\[9\] net844 net828 total_design.core.regFile.register\[1\]\[9\]
+ _02568_ vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_116_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06850__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload145 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 clkload145/Y sky130_fd_sc_hd__inv_8
XANTENNA__10715__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload156 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 clkload156/Y sky130_fd_sc_hd__inv_8
XFILLER_0_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload167 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 clkload167/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_168_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload178 clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 clkload178/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_105_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06602__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap999 net1000 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_1
X_08972_ net473 _02666_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__or2_1
XANTENNA__09364__X _04604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07923_ total_design.core.regFile.register\[15\]\[27\] net847 net820 total_design.core.regFile.register\[17\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__a22o_1
Xhold18 total_design.core.data_mem.data_read_adr_reg\[5\] vssd1 vssd1 vccd1 vccd1
+ net1334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 total_design.core.data_mem.data_read_adr_reg\[11\] vssd1 vssd1 vccd1 vccd1
+ net1345 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11546__S net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout197_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10450__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07854_ total_design.core.regFile.register\[29\]\[25\] net656 net567 total_design.core.regFile.register\[12\]\[25\]
+ _03356_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__a221o_1
X_06805_ total_design.core.regFile.register\[14\]\[5\] net626 net617 total_design.core.regFile.register\[10\]\[5\]
+ _02364_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07785_ total_design.core.regFile.register\[1\]\[24\] net828 net787 total_design.core.regFile.register\[13\]\[24\]
+ _03290_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__a221o_1
X_09524_ net903 _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__nor2_1
X_06736_ total_design.core.regFile.register\[10\]\[4\] net834 net763 total_design.core.regFile.register\[6\]\[4\]
+ _02299_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a221o_1
X_09455_ _04644_ _04690_ net461 vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06667_ net554 total_design.core.ctrl.imm_32\[2\] vssd1 vssd1 vccd1 vccd1 _02235_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout152_X net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout629_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ _03760_ _03761_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__or2_1
X_09386_ net314 _04432_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__nor2_1
XANTENNA__07881__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06598_ total_design.core.regFile.register\[18\]\[1\] net746 net737 net731 vssd1
+ vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08337_ total_design.core.data_mem.data_write_adr_reg\[26\] net546 net538 total_design.core.data_mem.data_read_adr_reg\[26\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08268_ net1391 net558 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[18\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_117_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07633__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07219_ total_design.core.regFile.register\[23\]\[13\] net681 net569 total_design.core.regFile.register\[17\]\[13\]
+ _02753_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__a221o_1
X_08199_ _03652_ _03653_ _03655_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__or3_1
X_10230_ net285 total_design.core.regFile.register\[15\]\[0\] net500 vssd1 vssd1 vccd1
+ vccd1 _00519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10161_ net275 net2084 net396 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1005 net1006 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09274__X _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_58_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1016 net1018 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1027 net1059 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__clkbuf_4
Xfanout1038 net1045 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10092_ net257 net2478 net403 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13882__D total_design.core.ctrl.imm_32\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11456__S net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1049 net1051 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13920_ clknet_leaf_82_clk _01100_ net1241 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10360__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13851_ clknet_leaf_52_clk _01059_ net1094 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12802_ clknet_leaf_126_clk _00269_ net1192 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13782_ clknet_leaf_50_clk total_design.core.data_mem.stored_data_adr\[25\] net1100
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[25\] sky130_fd_sc_hd__dfrtp_1
X_10994_ net520 _05252_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__nand2_2
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11653__A0 _05477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ clknet_leaf_9_clk _00200_ net1019 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06285__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12664_ clknet_leaf_134_clk _00131_ net1189 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14403_ clknet_leaf_47_clk net1876 net1097 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11615_ _05633_ net1768 net139 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12595_ clknet_leaf_179_clk _00062_ net1034 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14334_ clknet_leaf_52_clk _01495_ net1094 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[25\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07085__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11546_ net1617 _05643_ net146 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14265_ clknet_leaf_66_clk _01444_ net1122 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11477_ net1578 _05612_ net153 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__mux2_1
XANTENNA__10535__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13216_ clknet_leaf_193_clk _00683_ net1012 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10428_ net284 net2825 net381 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14196_ clknet_leaf_79_clk _01376_ net1221 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_164_Right_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13147_ clknet_leaf_144_clk _00614_ net1174 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ net167 total_design.core.regFile.register\[12\]\[30\] net490 vssd1 vssd1
+ vccd1 vccd1 _00645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13078_ clknet_leaf_155_clk _00545_ net1137 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13792__D total_design.core.data_mem.data_cpu_i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12029_ _05883_ _05885_ _05887_ _05889_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__or4_1
XANTENNA__10270__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07145__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__A0 total_design.core.math.pc_val\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06899__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ _03084_ _03064_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11644__A0 _05648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06521_ total_design.core.regFile.register\[3\]\[0\] net743 net737 net733 vssd1 vssd1
+ vccd1 vccd1 _02095_ sky130_fd_sc_hd__and4_1
XANTENNA__08805__A2_N _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09240_ _04216_ _04484_ net317 vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06452_ net973 _02025_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__nor2_1
XANTENNA__07863__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09171_ _04418_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__inv_2
X_06383_ net927 net911 net946 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__and3_4
XFILLER_0_44_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08122_ total_design.core.regFile.register\[31\]\[31\] net832 net777 total_design.core.regFile.register\[22\]\[31\]
+ _03613_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__a221o_1
XANTENNA__07615__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08812__A1 _02367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14522__1294 vssd1 vssd1 vccd1 vccd1 net1294 _14522__1294/LO sky130_fd_sc_hd__conb_1
X_08053_ total_design.core.regFile.register\[19\]\[29\] net640 _03547_ net686 vssd1
+ vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06823__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10445__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07004_ total_design.core.regFile.register\[22\]\[9\] net676 net614 total_design.core.regFile.register\[11\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11487__D _05479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08040__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1021_A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1119_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ _02188_ net703 _04207_ net533 vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__a211o_1
XANTENNA__06511__X _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout481_A _05011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ total_design.core.regFile.register\[22\]\[26\] net675 net667 total_design.core.regFile.register\[13\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__a22o_1
XANTENNA__10180__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08886_ net470 _02515_ _04139_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_99_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11883__A0 total_design.core.math.pc_val\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06597__C net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07000__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ total_design.core.regFile.register\[3\]\[25\] net867 net851 total_design.core.regFile.register\[9\]\[25\]
+ _03340_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__a221o_1
XFILLER_0_169_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07768_ _03273_ _03274_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__nand2b_1
XANTENNA__06894__A _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11635__A0 _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09507_ net207 net2491 net453 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__mux2_1
X_06719_ total_design.core.regFile.register\[18\]\[3\] net608 net589 total_design.core.regFile.register\[1\]\[3\]
+ _02268_ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07839__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ total_design.core.regFile.register\[20\]\[22\] net671 net571 total_design.core.regFile.register\[17\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09438_ _04663_ _04665_ _04674_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__or3b_1
XANTENNA__07854__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09369_ total_design.core.math.pc_val\[14\] _04583_ vssd1 vssd1 vccd1 vccd1 _04609_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_35_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11400_ net513 _05608_ _05656_ _05658_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12060__B1 _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12380_ _01639_ _01640_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__nand2_1
XANTENNA__07606__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08803__A1 total_design.core.data_mem.data_cpu_i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13877__D total_design.core.ctrl.imm_32\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11331_ _05530_ _05537_ _05448_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06814__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ clknet_leaf_87_clk _01230_ net1248 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11262_ _05514_ _05520_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13001_ clknet_leaf_16_clk _00468_ net1023 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10213_ _04759_ net2794 net391 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11193_ net513 _05271_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__nand2_1
XANTENNA__08031__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10144_ net193 net2255 net399 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__mux2_1
XANTENNA__06421__X _01997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10090__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10075_ net203 net2335 net407 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__mux2_1
X_13903_ clknet_leaf_84_clk _01083_ net1245 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11981__Y _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13834_ clknet_leaf_63_clk _01042_ net1122 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11626__A0 _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09180__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13765_ clknet_leaf_59_clk total_design.core.data_mem.stored_data_adr\[8\] net1126
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10977_ _05215_ _05231_ _05233_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08098__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12716_ clknet_leaf_167_clk _00183_ net1156 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13696_ clknet_leaf_40_clk total_design.core.data_mem.stored_read_data\[3\] net1091
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12647_ clknet_leaf_18_clk _00114_ net1047 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07058__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08083__X total_design.core.data_mem.data_cpu_i\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12578_ clknet_leaf_126_clk _00045_ net1193 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06805__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14317_ clknet_leaf_66_clk _01478_ net1123 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11529_ net1556 _05663_ net148 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10265__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold307 total_design.lcd_display.row_1\[88\] vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08243__B net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold318 total_design.lcd_display.row_2\[95\] vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold329 total_design.lcd_display.row_2\[49\] vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08007__C1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14248_ clknet_leaf_109_clk _01428_ net1231 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11885__A total_design.core.math.pc_val\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14179_ clknet_leaf_79_clk net1708 net1218 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08022__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout809 _01972_ vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__buf_4
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08740_ _03234_ _03282_ _03330_ _03995_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__and4_1
Xhold1007 total_design.core.regFile.register\[28\]\[2\] vssd1 vssd1 vccd1 vccd1 net2323
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 total_design.core.regFile.register\[24\]\[28\] vssd1 vssd1 vccd1 vccd1 net2334
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 total_design.core.regFile.register\[2\]\[28\] vssd1 vssd1 vccd1 vccd1 net2345
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08671_ total_design.lcd_display.cnt_500hz\[13\] total_design.lcd_display.cnt_500hz\[14\]
+ _03946_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__nand3_1
X_07622_ _03112_ _03132_ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11617__A0 _05651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07553_ total_design.core.regFile.register\[13\]\[19\] net787 net780 total_design.core.regFile.register\[27\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__a22o_1
XANTENNA__08089__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06504_ net744 net734 net728 vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07297__B1 _01959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07484_ total_design.core.regFile.register\[23\]\[18\] net678 net581 total_design.core.regFile.register\[6\]\[18\]
+ _03004_ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__a221o_1
XANTENNA__07836__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09223_ _04193_ _04463_ _04465_ _04468_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06435_ _02007_ _02008_ net690 _02010_ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__nand4_1
XFILLER_0_107_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1069_A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07049__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12042__B1 _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09154_ net257 net2233 net456 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__mux2_1
X_06366_ net966 net965 vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08105_ _03595_ _03597_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10175__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09085_ _04223_ _04227_ net464 vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06297_ _01808_ _01875_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09964__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08036_ total_design.core.regFile.register\[0\]\[29\] net873 _03531_ vssd1 vssd1
+ vccd1 vccd1 _03532_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold830 total_design.core.regFile.register\[26\]\[9\] vssd1 vssd1 vccd1 vccd1 net2146
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 total_design.core.regFile.register\[17\]\[22\] vssd1 vssd1 vccd1 vccd1 net2157
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold852 total_design.core.regFile.register\[6\]\[5\] vssd1 vssd1 vccd1 vccd1 net2168
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold863 total_design.core.regFile.register\[8\]\[27\] vssd1 vssd1 vccd1 vccd1 net2179
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 total_design.core.regFile.register\[23\]\[13\] vssd1 vssd1 vccd1 vccd1 net2190
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 total_design.core.regFile.register\[16\]\[11\] vssd1 vssd1 vccd1 vccd1 net2201
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 total_design.core.regFile.register\[21\]\[15\] vssd1 vssd1 vccd1 vccd1 net2212
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09265__A _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07221__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ net245 net1920 net415 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_A net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08600__C net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ _02337_ _04098_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__nand2_1
XANTENNA__06401__B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1530 total_design.core.regFile.register\[9\]\[10\] vssd1 vssd1 vccd1 vccd1 net2846
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09513__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1541 total_design.core.regFile.register\[29\]\[24\] vssd1 vssd1 vccd1 vccd1 net2857
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1552 total_design.core.regFile.register\[16\]\[23\] vssd1 vssd1 vccd1 vccd1 net2868
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ _01746_ _04097_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__or2_2
Xhold1563 total_design.core.regFile.register\[0\]\[18\] vssd1 vssd1 vccd1 vccd1 net2879
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10900_ _05132_ _05138_ _05158_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__a21o_1
X_11880_ total_design.core.math.pc_val\[0\] total_design.core.program_count.imm_val_reg\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11608__A0 _05609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10831_ _05076_ _05085_ _05079_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout916_X net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13550_ clknet_leaf_190_clk _01017_ net1034 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07288__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10762_ net2155 _05020_ _01775_ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07827__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12501_ net974 total_design.core.instr_mem.instruction_i\[14\] vssd1 vssd1 vccd1
+ vccd1 _01705_ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13481_ clknet_leaf_17_clk _00948_ net1046 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10874__A total_design.core.data_bus_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10693_ net247 net1903 net357 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__mux2_1
XANTENNA__08790__A_N total_design.core.data_mem.data_cpu_i\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12432_ net1895 net245 net344 vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__mux2_1
XANTENNA__12033__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06416__X _01992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12363_ _01613_ _01615_ _01616_ _01624_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__a211o_1
XANTENNA__10085__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14102_ clknet_leaf_101_clk _01282_ net1237 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11314_ net294 _05572_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_130_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09874__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11976__Y _05838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07460__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12294_ total_design.core.math.pc_val\[17\] total_design.core.program_count.imm_val_reg\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14033_ clknet_leaf_96_clk _01213_ net1253 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_11245_ _05399_ _05407_ _05500_ _05501_ _05502_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08004__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ _05422_ _05423_ _05429_ _05433_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__a31oi_1
XANTENNA__06566__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10127_ net274 net2746 net401 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10058_ net282 net2183 net406 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__mux2_1
XANTENNA__07515__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11644__S net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14521__1293 vssd1 vssd1 vccd1 vccd1 net1293 _14521__1293/LO sky130_fd_sc_hd__conb_1
XFILLER_0_54_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_106_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13817_ clknet_leaf_71_clk total_design.core.data_mem.data_cpu_i\[26\] net1206 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[26\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10120__Y _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11075__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07279__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13748_ clknet_leaf_72_clk total_design.core.data_mem.stored_write_data\[23\] net1220
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_57_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13679_ clknet_leaf_49_clk total_design.core.data_mem.data_read_adr_i\[19\] net1101
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[19\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06220_ total_design.core.instr_mem.instruction_adr_i\[8\] total_design.core.instr_mem.instruction_adr_stored\[8\]
+ net984 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__mux2_1
XANTENNA__12024__B1 _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06326__X _01905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06151_ net35 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09784__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold104 total_design.core.data_mem.data_bus_i_reg\[20\] vssd1 vssd1 vccd1 vccd1 net1420
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 total_design.core.instr_mem.instruction_adr_stored\[7\] vssd1 vssd1 vccd1
+ vccd1 net1431 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07451__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold126 total_design.core.data_mem.data_bus_i_reg\[21\] vssd1 vssd1 vccd1 vccd1 net1442
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold137 total_design.core.data_mem.data_bus_i_reg\[28\] vssd1 vssd1 vccd1 vccd1 net1453
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 total_design.core.data_mem.data_read_adr_reg2\[5\] vssd1 vssd1 vccd1 vccd1
+ net1464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold159 total_design.core.math.pc_val\[8\] vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ net181 net2519 net427 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10723__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout606 net607 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_4
X_09841_ net186 net2130 net436 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout617 net618 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout628 net631 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_8
Xfanout639 _02060_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09772_ net189 net2857 net444 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__mux2_1
X_06984_ total_design.core.regFile.register\[0\]\[8\] net876 _02520_ _02534_ vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[8\] sky130_fd_sc_hd__o22a_4
X_08723_ net115 net114 net112 net113 vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__nand4b_1
XPHY_EDGE_ROW_13_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout277_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11554__S net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08654_ total_design.lcd_display.cnt_500hz\[7\] total_design.lcd_display.cnt_500hz\[6\]
+ _03933_ total_design.lcd_display.cnt_500hz\[8\] vssd1 vssd1 vccd1 vccd1 _03938_
+ sky130_fd_sc_hd__a31o_1
X_07605_ total_design.core.regFile.register\[28\]\[20\] net853 net819 total_design.core.regFile.register\[17\]\[20\]
+ _03118_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08585_ _03822_ net880 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout444_A _04969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07536_ total_design.core.regFile.register\[22\]\[19\] net675 net617 total_design.core.regFile.register\[10\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__a22o_1
XANTENNA__09959__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06594__D net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07809__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07467_ _02969_ _02989_ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout611_A _02072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09206_ net265 net2288 net454 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__mux2_1
XANTENNA__12015__B1 _05839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06418_ net966 _01739_ net918 _01936_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__and4_4
XANTENNA__07690__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07398_ total_design.core.regFile.register\[2\]\[16\] net785 _02922_ _02924_ vssd1
+ vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__a211o_1
XFILLER_0_161_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11369__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09137_ net322 _04252_ _04385_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__o21ai_1
X_06349_ net951 net950 total_design.core.ctrl.instruction\[24\] net952 vssd1 vssd1
+ vccd1 vccd1 _01925_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ net705 _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__nor2_1
XANTENNA__07442__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout980_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06796__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ total_design.core.regFile.register\[19\]\[29\] net823 net767 total_design.core.regFile.register\[7\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__a22o_1
XANTENNA__10633__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10329__A0 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 total_design.core.regFile.register\[1\]\[15\] vssd1 vssd1 vccd1 vccd1 net1976
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold671 total_design.core.regFile.register\[30\]\[21\] vssd1 vssd1 vccd1 vccd1 net1987
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11030_ net351 _05055_ _05221_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__and3_1
Xhold682 total_design.core.regFile.register\[28\]\[15\] vssd1 vssd1 vccd1 vccd1 net1998
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 total_design.core.regFile.register\[26\]\[23\] vssd1 vssd1 vccd1 vccd1 net2009
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout866_X net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09723__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ clknet_leaf_157_clk _00448_ net1141 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11464__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09498__B2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1360 total_design.core.regFile.register\[9\]\[11\] vssd1 vssd1 vccd1 vccd1 net2676
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1371 total_design.core.regFile.register\[8\]\[10\] vssd1 vssd1 vccd1 vccd1 net2687
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11932_ total_design.keypad0.key_out\[12\] net529 _05797_ total_design.keypad0.key_out\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1382 total_design.core.regFile.register\[10\]\[0\] vssd1 vssd1 vccd1 vccd1 net2698
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1393 total_design.core.regFile.register\[21\]\[18\] vssd1 vssd1 vccd1 vccd1 net2709
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11863_ total_design.lcd_display.currentState\[2\] _05722_ vssd1 vssd1 vccd1 vccd1
+ _05747_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13602_ clknet_leaf_60_clk net1328 net1132 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10814_ _05061_ _05069_ _05070_ _05071_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__a31o_1
XANTENNA__09869__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11794_ net1781 net954 _05699_ _01791_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10745_ net2874 net353 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_60_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13533_ clknet_leaf_14_clk _01000_ net1026 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12006__B1 _05839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07681__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13464_ clknet_leaf_136_clk _00931_ net1181 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10676_ net214 net2388 net361 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12415_ total_design.core.math.pc_val\[30\] net989 vssd1 vssd1 vccd1 vccd1 _01672_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_91_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13395_ clknet_leaf_178_clk _00862_ net1035 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10568__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12346_ net990 _04779_ _01610_ net894 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__o211a_1
XANTENNA__07433__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11639__S net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12277_ _06113_ _06114_ _06116_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__or3_1
XANTENNA__10543__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14016_ clknet_leaf_111_clk _01196_ net1227 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_11228_ _05486_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__inv_2
XANTENNA_output73_A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11159_ _05414_ _05415_ _05417_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_147_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08948__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06711__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08370_ _03726_ _03727_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07321_ total_design.core.regFile.register\[18\]\[15\] net610 net572 total_design.core.regFile.register\[17\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10718__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09661__A1 total_design.core.ctrl.instruction\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09661__B2 total_design.core.data_cpu_o\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07252_ _02778_ _02783_ _02785_ _02787_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__or4_1
XFILLER_0_144_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06203_ total_design.core.data_adr_o\[15\] _01781_ net963 vssd1 vssd1 vccd1 vccd1
+ _01782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07183_ total_design.core.regFile.register\[26\]\[12\] net870 net764 total_design.core.regFile.register\[6\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10961__B net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11549__S net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10453__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09527__B _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout403 net405 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09716__A2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06232__A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout414 _04983_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_6
Xfanout425 _04979_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_8
Xfanout436 net437 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout394_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09824_ net261 net2260 net437 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__mux2_1
Xfanout447 _04189_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_2
Xfanout469 net470 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_2
X_09755_ net266 net2396 net443 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__mux2_1
X_06967_ total_design.core.regFile.register\[15\]\[8\] net848 net844 total_design.core.regFile.register\[25\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout659_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06950__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ net2583 _03952_ vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__xor2_1
X_09686_ _03487_ _03506_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__and2b_1
XANTENNA__08159__A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06898_ total_design.core.regFile.register\[13\]\[7\] net666 net663 total_design.core.regFile.register\[9\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a22o_1
X_08637_ total_design.lcd_display.cnt_500hz\[3\] total_design.lcd_display.cnt_500hz\[4\]
+ _03921_ _03925_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__and4b_1
XFILLER_0_139_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ total_design.data_in_BUS\[23\] net340 net719 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[23\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_30_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07519_ _02949_ _02991_ _02990_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_147_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08499_ _03845_ _03849_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__or2_1
XANTENNA__10628__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout614_X net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10530_ net269 net2072 net373 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_1054 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10461_ net284 net2137 net380 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__mux2_1
X_12200_ _04424_ _05757_ _05760_ _06048_ net526 vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_0_0_clk_X clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13180_ clknet_leaf_10_clk _00647_ net1021 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14520__1292 vssd1 vssd1 vccd1 vccd1 net1292 _14520__1292/LO sky130_fd_sc_hd__conb_1
XFILLER_0_33_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10392_ net168 net1962 net487 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout983_X net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06769__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11762__A2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11459__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ total_design.lcd_display.row_1\[46\] _05821_ _05829_ total_design.lcd_display.row_1\[110\]
+ _05986_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__a221o_1
XANTENNA__10363__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12062_ total_design.lcd_display.row_1\[19\] _05826_ _05844_ total_design.lcd_display.row_2\[43\]
+ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__a22o_1
Xhold490 total_design.lcd_display.row_2\[72\] vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11013_ net520 _05271_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__nand2_2
XANTENNA__06499__D net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout970 total_design.core.ctrl.instruction\[13\] vssd1 vssd1 vccd1 vccd1 net970
+ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07525__X total_design.core.ctrl.imm_32\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07194__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout981 net982 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_4
Xfanout992 net996 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06288__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12964_ clknet_leaf_105_clk _00431_ net1233 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1190 total_design.core.regFile.register\[28\]\[7\] vssd1 vssd1 vccd1 vccd1 net2506
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_103_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09740__X _04963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11915_ _05777_ _05791_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ clknet_leaf_183_clk _00362_ net1039 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _03928_ _05732_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11777_ net1740 net953 _05694_ _01830_ vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__a22o_1
X_14565_ net37 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10538__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11450__A1 _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10728_ total_design.core.regFile.register\[0\]\[3\] net355 vssd1 vssd1 vccd1 vccd1
+ _01002_ sky130_fd_sc_hd__and2_1
XANTENNA__07654__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13516_ clknet_leaf_164_clk _00983_ net1158 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07420__B total_design.core.ctrl.instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_125_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14496_ clknet_leaf_33_clk _01563_ net1072 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_24_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13447_ clknet_leaf_176_clk _00914_ net1048 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10659_ net286 net2507 net364 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__mux2_1
Xclkload13 clknet_leaf_198_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_35_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload24 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload24/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__06209__A1 _01771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload35 clknet_leaf_189_clk vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07406__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload46 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_51_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13378_ clknet_leaf_129_clk _00845_ net1193 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload57 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__inv_8
XANTENNA__13795__D total_design.core.data_mem.data_cpu_i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkload68 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__inv_8
XFILLER_0_51_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload79 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_77_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12329_ total_design.core.math.pc_val\[20\] total_design.core.program_count.imm_val_reg\[20\]
+ _01591_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__a21boi_1
XANTENNA__10273__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07148__A _02666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07870_ _03371_ _03372_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__nand2b_2
XANTENNA__07185__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06821_ total_design.core.regFile.register\[12\]\[5\] net773 net771 total_design.core.regFile.register\[28\]\[5\]
+ _02380_ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a221o_1
X_09540_ net320 _04599_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__nor2_1
X_06752_ total_design.core.ctrl.instruction\[24\] _02311_ _02314_ vssd1 vssd1 vccd1
+ vccd1 total_design.core.ctrl.imm_32\[4\] sky130_fd_sc_hd__a21o_1
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09471_ _03088_ net537 _04188_ _03087_ _04705_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__a221o_1
X_06683_ total_design.core.regFile.register\[23\]\[3\] net811 _02249_ vssd1 vssd1
+ vccd1 vccd1 _02250_ sky130_fd_sc_hd__a21o_1
X_14544__1316 vssd1 vssd1 vccd1 vccd1 net1316 _14544__1316/LO sky130_fd_sc_hd__conb_1
X_08422_ _03773_ _03776_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11404__Y _05663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08353_ _03710_ _03712_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10448__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14203__RESET_B net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07304_ _02827_ _02829_ _02831_ _02836_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__or4_1
XANTENNA__11441__A1 _05652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08284_ _03658_ net561 vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__nor2_2
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload7 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_8
XFILLER_0_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06999__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11992__A2 _05832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07235_ total_design.core.regFile.register\[0\]\[13\] net873 vssd1 vssd1 vccd1 vccd1
+ _02771_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout407_A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1149_A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07166_ total_design.core.regFile.register\[30\]\[12\] net660 net582 total_design.core.regFile.register\[6\]\[12\]
+ _02704_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__a221o_1
XANTENNA__11744__A2 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10183__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08070__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07097_ net751 _02640_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[10\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09972__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout200 _04783_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_2
Xfanout1209 net1210 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__clkbuf_4
Xfanout211 _04721_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout776_A _01990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout222 net223 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__buf_1
Xfanout233 net235 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
Xfanout244 net245 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_2
Xfanout255 net256 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07176__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout266 _04452_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_2
X_09807_ net181 total_design.core.regFile.register\[28\]\[26\] net439 vssd1 vssd1
+ vccd1 vccd1 _00129_ sky130_fd_sc_hd__mux2_1
Xfanout277 net279 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__buf_1
XANTENNA_fanout943_A _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07999_ total_design.core.regFile.register\[14\]\[28\] net625 net578 total_design.core.regFile.register\[27\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06923__A2 _01949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09738_ _04193_ _04960_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ _03512_ net704 _04894_ net535 vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11700_ net4 net935 net878 net1509 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__o22a_1
XFILLER_0_167_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12209__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06687__B2 _01932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12680_ clknet_leaf_173_clk _00147_ net1055 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11631_ _05670_ net1776 net136 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__mux2_1
XANTENNA__10358__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11432__A1 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14350_ clknet_leaf_45_clk _00037_ net1086 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11562_ _05663_ net1784 net142 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__mux2_1
XANTENNA__07636__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10513_ net209 net2186 net482 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__mux2_1
X_13301_ clknet_leaf_161_clk _00768_ net1143 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14281_ net987 _01457_ net1082 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11493_ net1636 _05626_ net152 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13232_ clknet_leaf_182_clk _00699_ net1038 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09389__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10444_ net220 net1922 net382 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ clknet_leaf_107_clk _00630_ net1224 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10375_ net229 net2064 net484 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12114_ _05813_ _05825_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__nor2_1
XANTENNA__11984__Y _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13094_ clknet_leaf_195_clk _00561_ net1008 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11499__A1 _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12045_ total_design.lcd_display.row_2\[66\] _05819_ _05853_ total_design.lcd_display.row_2\[114\]
+ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07167__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09183__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06914__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13996_ clknet_leaf_99_clk _01176_ net1241 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12947_ clknet_leaf_190_clk _00414_ net1034 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07875__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12878_ clknet_leaf_187_clk _00345_ net1031 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10268__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11829_ total_design.lcd_display.cnt_20ms\[15\] _05715_ total_design.lcd_display.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11423__A1 _05626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10226__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07627__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14548_ net1268 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_126_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14479_ clknet_leaf_36_clk _01546_ net1072 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkload102 clknet_leaf_156_clk vssd1 vssd1 vccd1 vccd1 clkload102/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload113 clknet_leaf_163_clk vssd1 vssd1 vccd1 vccd1 clkload113/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07020_ total_design.core.regFile.register\[8\]\[9\] net804 net780 total_design.core.regFile.register\[27\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload124 clknet_leaf_139_clk vssd1 vssd1 vccd1 vccd1 clkload124/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_116_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload135 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 clkload135/Y sky130_fd_sc_hd__clkinv_2
Xclkload146 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 clkload146/X sky130_fd_sc_hd__clkbuf_8
Xclkload157 clknet_leaf_80_clk vssd1 vssd1 vccd1 vccd1 clkload157/Y sky130_fd_sc_hd__inv_6
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_168_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload168 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 clkload168/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_168_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload179 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 clkload179/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__08052__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09792__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08971_ _04220_ _04223_ net464 vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__mux2_1
X_07922_ total_design.core.regFile.register\[14\]\[27\] net862 net835 total_design.core.regFile.register\[10\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__a22o_1
Xhold19 total_design.core.data_mem.data_read_adr_reg\[31\] vssd1 vssd1 vccd1 vccd1
+ net1335 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12151__A2 _05834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ total_design.core.regFile.register\[26\]\[25\] net646 net574 total_design.core.regFile.register\[24\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06905__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14500__Q total_design.core.ctrl.instruction\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_06804_ total_design.core.regFile.register\[27\]\[5\] net579 net564 total_design.core.regFile.register\[3\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__a22o_1
X_07784_ total_design.core.regFile.register\[8\]\[24\] net803 net760 total_design.core.regFile.register\[21\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09523_ total_design.core.math.pc_val\[21\] _04735_ vssd1 vssd1 vccd1 vccd1 _04756_
+ sky130_fd_sc_hd__xnor2_1
X_06735_ total_design.core.regFile.register\[25\]\[4\] net842 net802 total_design.core.regFile.register\[8\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__a22o_1
XANTENNA__11562__S net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_A _05017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06669__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ _02969_ net308 net334 vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__mux2_1
X_06666_ net333 vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07330__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08405_ _03758_ _03759_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10178__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09385_ _04443_ _04623_ net319 vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__mux2_1
XANTENNA__09607__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06597_ total_design.core.regFile.register\[19\]\[1\] net746 net737 net732 vssd1
+ vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__and4_1
XANTENNA__08156__B _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1266_A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ net1493 net938 _03702_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[25\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09967__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09083__A2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08267_ net1371 net557 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[17\]
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout312_X net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_140_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_140_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ total_design.core.regFile.register\[2\]\[13\] net636 net620 total_design.core.regFile.register\[4\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__a22o_1
XANTENNA__06841__A1 total_design.core.ctrl.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_61_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08172__A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08198_ total_design.core.data_mem.data_write_adr_reg\[13\] total_design.core.data_mem.data_write_adr_reg\[12\]
+ total_design.core.data_mem.data_write_adr_reg\[15\] total_design.core.data_mem.data_write_adr_reg\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout893_A _02022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08603__C net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07149_ _02666_ _02688_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__nand2_1
XANTENNA__08043__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1221_X net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07397__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10160_ net258 net2861 net396 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 net1027 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ net280 total_design.core.regFile.register\[19\]\[4\] net402 vssd1 vssd1 vccd1
+ vccd1 _00395_ sky130_fd_sc_hd__mux2_1
Xfanout1017 net1018 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10641__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1028 net1029 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1039 net1045 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12142__A2 _05814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07516__A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06420__A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout946_X net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13850_ clknet_leaf_52_clk _01058_ net1094 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07235__B net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14196__RESET_B net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12801_ clknet_leaf_122_clk _00268_ net1167 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13781_ clknet_leaf_48_clk total_design.core.data_mem.stored_data_adr\[24\] net1099
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[24\] sky130_fd_sc_hd__dfrtp_1
X_10993_ total_design.core.data_bus_o\[2\] net696 vssd1 vssd1 vccd1 vccd1 _05252_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_172_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11472__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07857__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12732_ clknet_leaf_10_clk _00199_ net1019 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06419__X _01995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07321__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12663_ clknet_leaf_163_clk _00130_ net1166 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10088__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14402_ clknet_leaf_50_clk net1382 net1097 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09877__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11614_ _05646_ net1644 net140 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__mux2_1
XANTENNA__11979__Y _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_187_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12594_ clknet_leaf_146_clk _00061_ net1177 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14333_ clknet_leaf_52_clk _01494_ net1093 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[24\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_137_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11545_ net1788 _05648_ net145 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_131_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09178__A _04121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11476_ net1539 _05609_ net155 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__mux2_1
X_14264_ clknet_leaf_102_clk _01443_ net1239 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.currentState\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13215_ clknet_leaf_155_clk _00682_ net1137 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10427_ _04976_ net532 vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14195_ clknet_leaf_111_clk _01375_ net1208 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_150_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14543__1315 vssd1 vssd1 vccd1 vccd1 net1315 _14543__1315/LO sky130_fd_sc_hd__conb_1
XANTENNA__07388__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09782__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10358_ net171 net2712 net488 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__mux2_1
X_13146_ clknet_leaf_125_clk _00613_ net1188 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08810__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11647__S net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10551__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13077_ clknet_leaf_159_clk _00544_ net1143 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_163_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ net181 net1992 net498 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_125_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12133__A2 _05834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12028_ total_design.lcd_display.row_1\[73\] _05816_ _05873_ _05888_ vssd1 vssd1
+ vccd1 vccd1 _05889_ sky130_fd_sc_hd__a211o_1
XANTENNA__11219__Y _05478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06330__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_198_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_198_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06348__B1 _01915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_2__f_clk_X clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09641__A _03467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07560__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13979_ clknet_leaf_93_clk _01159_ net1255 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06520_ net740 net737 net732 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__and3_1
XANTENNA__07848__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06451_ total_design.core.ctrl.instruction\[4\] net972 _01915_ vssd1 vssd1 vccd1
+ vccd1 _02025_ sky130_fd_sc_hd__or3_2
XFILLER_0_75_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09787__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09170_ _04288_ _04417_ net327 vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_118_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06382_ net922 net917 net913 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08121_ total_design.core.regFile.register\[29\]\[31\] net799 net784 total_design.core.regFile.register\[2\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_122_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08812__A2 _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08052_ total_design.core.regFile.register\[8\]\[29\] net593 net585 total_design.core.regFile.register\[28\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__a22o_1
X_07003_ total_design.core.regFile.register\[10\]\[9\] net618 _02550_ vssd1 vssd1
+ vccd1 vccd1 _02551_ sky130_fd_sc_hd__a21o_1
XANTENNA__08025__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07379__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11580__A0 _05645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11557__S net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10461__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ _04205_ _04206_ net703 vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1014_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12124__A2 _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ total_design.core.regFile.register\[1\]\[26\] net590 net586 total_design.core.regFile.register\[28\]\[26\]
+ _03405_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_189_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_189_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08885_ net334 _02564_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__nor2_1
X_07836_ total_design.core.regFile.register\[19\]\[25\] net824 net807 total_design.core.regFile.register\[5\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__a22o_1
XANTENNA__07551__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ net554 total_design.core.data_mem.data_cpu_i\[23\] total_design.core.ctrl.imm_32\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout641_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09506_ _04734_ _04739_ net506 vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__o21a_2
XFILLER_0_149_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06718_ total_design.core.regFile.register\[19\]\[3\] net641 net597 total_design.core.regFile.register\[21\]\[3\]
+ _02272_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__a221o_1
XANTENNA__07839__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08167__A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07698_ net553 _03206_ _03179_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07303__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06649_ total_design.core.regFile.register\[23\]\[2\] net678 net608 total_design.core.regFile.register\[18\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__a22o_1
X_09437_ _02991_ net447 _04216_ _04664_ _04673_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__o221a_1
XFILLER_0_164_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout906_A _02014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ _04595_ _04607_ net449 vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_43_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08319_ total_design.core.data_mem.data_write_adr_reg\[17\] net547 net539 total_design.core.data_mem.data_read_adr_reg\[17\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__a221o_1
X_09299_ total_design.core.data_cpu_o\[11\] net757 _04541_ net906 _04538_ vssd1 vssd1
+ vccd1 vccd1 _04542_ sky130_fd_sc_hd__a221o_1
XANTENNA__10636__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_113_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_145_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08803__A2 _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13__f_clk_X clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11330_ _05576_ _05588_ _05538_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__or3b_1
X_11261_ _05427_ _05429_ _05516_ _05518_ _05519_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__a32o_2
XTAP_TAPCELL_ROW_132_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10212_ net208 net2195 net389 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__mux2_1
X_13000_ clknet_leaf_172_clk _00467_ net1056 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07224__D1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09726__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ net513 _05271_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11467__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ net197 net2692 net400 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__mux2_1
XANTENNA__10371__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07790__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_A gpio_in[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ net207 net1938 net406 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13902_ clknet_leaf_111_clk _01082_ net1209 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07542__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13833_ clknet_leaf_59_clk _01041_ net1127 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13764_ clknet_leaf_60_clk total_design.core.data_mem.stored_data_adr\[7\] net1132
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10976_ _05231_ _05233_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_139_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12715_ clknet_leaf_127_clk _00182_ net1191 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13695_ clknet_leaf_40_clk total_design.core.data_mem.stored_read_data\[2\] net1093
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12646_ clknet_leaf_200_clk _00113_ net1002 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10546__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_104_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12577_ clknet_leaf_121_clk _00044_ net1170 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09452__C1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14316_ clknet_leaf_63_clk _01477_ net1124 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_123_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11528_ net1564 _05627_ net147 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold308 total_design.lcd_display.row_2\[111\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold319 total_design.data_in_BUS\[27\] vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09204__C1 _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14247_ clknet_leaf_108_clk _01427_ net1231 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11459_ net1536 _05624_ net154 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11562__A0 _05663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ clknet_leaf_114_clk _01358_ net1208 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_2
XANTENNA__10281__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13129_ clknet_leaf_16_clk _00596_ net1023 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12106__A2 _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07781__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07156__A total_design.core.ctrl.instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1008 total_design.core.regFile.register\[16\]\[16\] vssd1 vssd1 vccd1 vccd1 net2324
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1019 total_design.core.regFile.register\[20\]\[21\] vssd1 vssd1 vccd1 vccd1 net2335
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08670_ total_design.lcd_display.cnt_500hz\[13\] total_design.lcd_display.cnt_500hz\[12\]
+ _03944_ total_design.lcd_display.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 _03948_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07533__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ _03112_ _03132_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__nand2_1
XANTENNA__06741__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07552_ total_design.core.regFile.register\[3\]\[19\] net867 _03068_ _03069_ vssd1
+ vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06503_ total_design.core.regFile.register\[31\]\[0\] net747 net733 net727 vssd1
+ vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__and4_1
X_07483_ total_design.core.regFile.register\[21\]\[18\] net597 net585 total_design.core.regFile.register\[28\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09222_ _02539_ net508 net298 _04466_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__o221ai_1
X_06434_ _01740_ _01993_ _01960_ _01946_ net874 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_174_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11412__Y _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09153_ net507 _04401_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06365_ net920 net948 net911 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__and3_4
XFILLER_0_17_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10456__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08797__A1 _02565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08104_ net553 total_design.core.data_mem.data_cpu_i\[30\] total_design.core.ctrl.imm_32\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09084_ _04258_ _04220_ net464 vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__mux2_1
XANTENNA__06235__A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06296_ net964 _01874_ _01873_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08035_ _03523_ _03525_ _03530_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold820 total_design.core.regFile.register\[15\]\[28\] vssd1 vssd1 vccd1 vccd1 net2136
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1131_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold831 total_design.core.regFile.register\[19\]\[21\] vssd1 vssd1 vccd1 vccd1 net2147
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1229_A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold842 total_design.core.regFile.register\[10\]\[27\] vssd1 vssd1 vccd1 vccd1 net2158
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 total_design.core.regFile.register\[18\]\[27\] vssd1 vssd1 vccd1 vccd1 net2169
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 total_design.core.regFile.register\[12\]\[19\] vssd1 vssd1 vccd1 vccd1 net2180
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 total_design.core.regFile.register\[23\]\[11\] vssd1 vssd1 vccd1 vccd1 net2191
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold886 total_design.data_in_BUS\[1\] vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10191__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold897 total_design.core.regFile.register\[23\]\[9\] vssd1 vssd1 vccd1 vccd1 net2213
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ net287 net1986 net414 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09980__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ _02338_ _04099_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06980__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout856_A _01947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06401__C net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1520 total_design.core.regFile.register\[13\]\[8\] vssd1 vssd1 vccd1 vccd1 net2836
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 total_design.core.regFile.register\[23\]\[30\] vssd1 vssd1 vccd1 vccd1 net2847
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 total_design.core.regFile.register\[11\]\[31\] vssd1 vssd1 vccd1 vccd1 net2858
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1553 total_design.core.regFile.register\[0\]\[27\] vssd1 vssd1 vccd1 vccd1 net2869
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08868_ _04118_ _04119_ _04114_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__or3b_4
Xhold1564 total_design.data_in_BUS\[11\] vssd1 vssd1 vccd1 vccd1 net2880 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07819_ _03303_ _03322_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__nor2_1
XANTENNA__06732__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08799_ _04052_ _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_28_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10830_ _05061_ _05087_ _05086_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542__1314 vssd1 vssd1 vccd1 vccd1 net1314 _14542__1314/LO sky130_fd_sc_hd__conb_1
XFILLER_0_165_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10761_ _01763_ _01772_ _05021_ total_design.core.data_access vssd1 vssd1 vccd1 vccd1
+ _01032_ sky130_fd_sc_hd__a22o_1
XANTENNA__12281__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_X net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout909_X net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12500_ net979 net970 net883 _01704_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13480_ clknet_leaf_24_clk _00947_ net1057 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10692_ net284 total_design.core.regFile.register\[1\]\[0\] net357 vssd1 vssd1 vccd1
+ vccd1 _00967_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12431_ total_design.core.regFile.register\[31\]\[0\] net284 net344 vssd1 vssd1 vccd1
+ vccd1 _01502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10366__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12362_ _01613_ _01616_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11792__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14101_ clknet_leaf_89_clk _01281_ net1258 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11313_ _05531_ _05568_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__xor2_1
X_12293_ _06122_ _06127_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__and2_1
X_11244_ _05501_ _05502_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__and2_1
X_14032_ clknet_leaf_110_clk _01212_ net1227 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09456__A _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ _05426_ _05429_ _05433_ _05424_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_101_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09890__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07763__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ net257 net2366 net400 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__mux2_1
XANTENNA__09743__X _04966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06971__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ net269 net2008 net407 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07515__A2 total_design.core.data_mem.data_cpu_i\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06723__B1 _02266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload0_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13816_ clknet_leaf_71_clk total_design.core.data_mem.data_cpu_i\[25\] net1205 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[25\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09268__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11075__A2 _05049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13747_ clknet_leaf_111_clk total_design.core.data_mem.stored_write_data\[22\] net1208
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[22\] sky130_fd_sc_hd__dfrtp_1
X_10959_ net521 _05184_ _05191_ _05187_ _05181_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__a32o_1
XANTENNA__11660__S net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13678_ clknet_leaf_49_clk total_design.core.data_mem.data_read_adr_i\[18\] net1101
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[18\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10276__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12629_ clknet_leaf_166_clk _00096_ net1157 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08254__B net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06150_ net2263 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold105 total_design.core.math.pc_val\[27\] vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 total_design.core.instr_mem.instruction_adr_stored\[14\] vssd1 vssd1 vccd1
+ vccd1 net1432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold127 total_design.core.instr_mem.instruction_adr_stored\[28\] vssd1 vssd1 vccd1
+ vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 total_design.core.data_mem.data_read_adr_reg2\[23\] vssd1 vssd1 vccd1 vccd1
+ net1454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 total_design.core.data_mem.data_read_adr_reg2\[3\] vssd1 vssd1 vccd1 vccd1
+ net1465 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12327__A2 _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09840_ net191 net2192 net436 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__mux2_1
Xfanout607 _02074_ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__buf_4
Xfanout618 net619 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_8
Xfanout629 net631 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07754__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09771_ net196 net2735 net442 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06983_ _02526_ _02528_ _02533_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__or3_1
XANTENNA__06962__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08722_ net115 net114 net112 net113 vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__and4b_1
XANTENNA__09813__B total_design.core.ctrl.instruction\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07506__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ net2864 _03936_ _03937_ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__o21a_1
XANTENNA__06714__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07604_ total_design.core.regFile.register\[14\]\[20\] net861 net850 total_design.core.regFile.register\[9\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08584_ _03796_ net880 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12263__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07535_ total_design.core.regFile.register\[11\]\[19\] net613 net586 total_design.core.regFile.register\[28\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1081_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11570__S net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout437_A _04973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1179_A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07466_ net551 net309 _02948_ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__o21a_1
XANTENNA__06517__X _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09205_ net452 _04451_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__nor2_2
X_06417_ _01738_ total_design.core.ctrl.instruction\[23\] net923 _01928_ vssd1 vssd1
+ vccd1 vccd1 _01993_ sky130_fd_sc_hd__or4_1
XFILLER_0_107_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10186__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07397_ total_design.core.regFile.register\[14\]\[16\] net862 net777 total_design.core.regFile.register\[22\]\[16\]
+ _02923_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout604_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08164__B _02492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09975__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06348_ _01917_ _01920_ _01915_ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__a21oi_4
X_09136_ net328 _04274_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08732__X total_design.lcd_display.lcd_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09067_ _02291_ _04317_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__xor2_1
X_06279_ net930 _01857_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1134_X net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08018_ total_design.core.regFile.register\[11\]\[29\] net794 net783 total_design.core.regFile.register\[2\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__a22o_1
XANTENNA__07993__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold650 total_design.core.regFile.register\[6\]\[26\] vssd1 vssd1 vccd1 vccd1 net1966
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout973_A total_design.core.ctrl.instruction\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout594_X net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 total_design.core.regFile.register\[20\]\[13\] vssd1 vssd1 vccd1 vccd1 net1977
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold672 total_design.core.regFile.register\[31\]\[9\] vssd1 vssd1 vccd1 vccd1 net1988
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold683 total_design.core.regFile.register\[31\]\[17\] vssd1 vssd1 vccd1 vccd1 net1999
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 total_design.core.regFile.register\[14\]\[28\] vssd1 vssd1 vccd1 vccd1 net2010
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07745__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ net213 net2878 net418 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06953__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_X net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ clknet_leaf_140_clk _00447_ net1182 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1350 total_design.core.regFile.register\[6\]\[21\] vssd1 vssd1 vccd1 vccd1 net2666
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1361 total_design.core.regFile.register\[5\]\[18\] vssd1 vssd1 vccd1 vccd1 net2677
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ total_design.keypad0.key_out\[11\] net529 net475 total_design.keypad0.key_out\[7\]
+ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__a22o_1
Xhold1372 total_design.core.regFile.register\[9\]\[14\] vssd1 vssd1 vccd1 vccd1 net2688
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06705__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1383 total_design.core.regFile.register\[11\]\[16\] vssd1 vssd1 vccd1 vccd1 net2699
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1394 total_design.core.regFile.register\[26\]\[7\] vssd1 vssd1 vccd1 vccd1 net2710
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11862_ total_design.lcd_display.currentState\[2\] _05745_ net709 vssd1 vssd1 vccd1
+ vccd1 _01440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13601_ clknet_leaf_61_clk net1334 net1129 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13533__RESET_B net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10813_ _05061_ _05069_ _05070_ _05071_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__a31oi_2
XANTENNA__12254__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ net1750 net955 net301 _01780_ vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__a22o_1
XANTENNA__11480__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13532_ clknet_leaf_28_clk _00999_ net1075 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_10744_ total_design.core.regFile.register\[0\]\[19\] net355 vssd1 vssd1 vccd1 vccd1
+ _01018_ sky130_fd_sc_hd__and2_1
XANTENNA__07130__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13463_ clknet_leaf_124_clk _00930_ net1186 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10096__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10675_ net222 net2132 net363 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__mux2_1
XANTENNA__09885__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12414_ total_design.core.math.pc_val\[29\] net524 _01665_ _01671_ vssd1 vssd1 vccd1
+ vccd1 _01499_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11987__Y _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13394_ clknet_leaf_139_clk _00861_ net1184 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06323__C_N _01900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12345_ _01597_ _01606_ _01607_ _01609_ vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08091__D1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07984__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12276_ total_design.core.math.pc_val\[15\] total_design.core.program_count.imm_val_reg\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__nor2_1
X_14015_ clknet_leaf_97_clk _01195_ net1244 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_11227_ _05386_ _05388_ _05483_ _05482_ _05372_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__a311o_1
XANTENNA__07736__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11158_ _05404_ _05416_ _05407_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_147_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11655__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10109_ net199 net2196 net403 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__mux2_1
X_11089_ _05346_ _05347_ net180 vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08146__C1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09125__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_159_Right_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08249__B _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12245__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10795__A total_design.core.data_bus_o\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07320_ total_design.core.regFile.register\[30\]\[15\] net661 net603 total_design.core.regFile.register\[31\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_173_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07121__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07251_ total_design.core.regFile.register\[13\]\[13\] net786 net779 total_design.core.regFile.register\[27\]\[13\]
+ _02786_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10008__A0 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06202_ total_design.core.instr_mem.instruction_adr_i\[15\] total_design.core.instr_mem.instruction_adr_stored\[15\]
+ net983 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09795__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07182_ total_design.core.regFile.register\[29\]\[12\] net798 net776 total_design.core.regFile.register\[22\]\[12\]
+ _02719_ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__a221o_1
XFILLER_0_170_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07975__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09177__B2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14541__1313 vssd1 vssd1 vccd1 vccd1 net1313 _14541__1313/LO sky130_fd_sc_hd__conb_1
Xfanout404 net405 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07188__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout415 _04983_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07727__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout426 net429 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_8
X_09823_ net267 net2632 net434 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__mux2_1
Xfanout437 _04973_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_8
Xfanout448 _04189_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__clkbuf_4
Xfanout459 net462 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_2
XANTENNA__06935__B1 _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11565__S net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__A_N _02818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ net273 net2575 net445 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06966_ total_design.core.regFile.register\[18\]\[8\] net858 net800 total_design.core.regFile.register\[29\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__a22o_1
X_08705_ _00029_ _00028_ _03970_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__or3_1
XANTENNA__12484__A1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09685_ net175 net2362 net455 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__mux2_1
X_06897_ total_design.core.regFile.register\[31\]\[7\] net601 net580 total_design.core.regFile.register\[27\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout554_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08159__B _02241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_93_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10495__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_169_Left_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08636_ total_design.lcd_display.cnt_500hz\[5\] total_design.lcd_display.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__nor2_1
XANTENNA__07360__B1 total_design.core.ctrl.imm_32\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12236__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ total_design.data_in_BUS\[22\] net341 net719 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[22\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_76_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1084_X net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout819_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07518_ _03036_ _03037_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__and2_2
XFILLER_0_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08498_ _03845_ _03849_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__nand2_1
XANTENNA__07112__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11995__B1 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08606__C net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07449_ total_design.core.regFile.register\[10\]\[17\] net834 net786 total_design.core.regFile.register\[13\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__a22o_1
XANTENNA__12997__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06407__B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ _04978_ net532 vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09404__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11747__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09119_ net298 _04357_ _04362_ net297 vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__o22a_1
XANTENNA__10644__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10391_ net169 net2817 net484 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12130_ total_design.lcd_display.row_1\[102\] _05810_ _05814_ total_design.lcd_display.row_1\[118\]
+ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06423__A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12061_ total_design.lcd_display.row_2\[91\] _05837_ _05841_ total_design.lcd_display.row_1\[11\]
+ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__a221o_1
Xhold480 total_design.data_in_BUS\[13\] vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold491 total_design.core.math.pc_val\[15\] vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ total_design.core.data_bus_o\[1\] net696 vssd1 vssd1 vccd1 vccd1 _05271_
+ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_53_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06926__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout960 _01911_ vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__buf_4
Xfanout971 net972 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__buf_2
Xfanout982 net985 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_4
Xfanout993 net996 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12963_ clknet_leaf_8_clk _00430_ net1016 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_84_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_142_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1180 total_design.core.regFile.register\[13\]\[23\] vssd1 vssd1 vccd1 vccd1 net2496
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08143__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1191 total_design.core.regFile.register\[2\]\[0\] vssd1 vssd1 vccd1 vccd1 net2507
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09340__A1 _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11914_ _03907_ _05773_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_142_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ clknet_leaf_167_clk _00361_ net1155 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11845_ total_design.lcd_display.currentState\[5\] _05731_ _05726_ vssd1 vssd1 vccd1
+ vccd1 _05732_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_157_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14564_ net36 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11776_ net1763 net954 _05699_ _01798_ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__a22o_1
XANTENNA__13699__Q total_design.core.data_cpu_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13515_ clknet_leaf_119_clk _00982_ net1171 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10727_ total_design.core.regFile.register\[0\]\[2\] net353 vssd1 vssd1 vccd1 vccd1
+ _01001_ sky130_fd_sc_hd__and2_1
X_14495_ clknet_leaf_27_clk _01562_ net1074 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08851__B1 _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13446_ clknet_leaf_199_clk _00913_ net1001 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10658_ _04989_ net532 vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__nand2_1
Xclkload14 clknet_leaf_199_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__inv_6
XFILLER_0_152_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload25 clknet_leaf_178_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_113_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload36 clknet_leaf_190_clk vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__10554__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13377_ clknet_leaf_118_clk _00844_ net1169 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload47 clknet_leaf_171_clk vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_140_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10589_ net170 net2725 net369 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__mux2_1
Xclkload58 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__inv_8
XFILLER_0_106_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload69 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__inv_6
XFILLER_0_24_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07957__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12328_ total_design.core.math.pc_val\[20\] net522 _01593_ _01594_ vssd1 vssd1 vccd1
+ vccd1 _01490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_149_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09159__A1 _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12259_ _06098_ _06099_ _06100_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__or3_1
XANTENNA__07709__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_166_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06620__X _02190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06917__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ total_design.core.regFile.register\[20\]\[5\] net817 _01969_ total_design.core.regFile.register\[4\]\[5\]
+ net693 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a221o_1
XANTENNA__07590__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06751_ total_design.core.ctrl.instruction\[11\] _01918_ net886 total_design.core.ctrl.instruction\[16\]
+ _02313_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_75_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08134__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09470_ _03084_ net505 vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__nor2_1
X_06682_ total_design.core.regFile.register\[20\]\[3\] net818 net775 total_design.core.regFile.register\[22\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a22o_1
XANTENNA_wire310_X net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07342__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08421_ _03753_ _03774_ _03775_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__or3_1
XANTENNA__06696__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11414__A _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08352_ total_design.data_from_keypad\[0\] _01888_ _03711_ vssd1 vssd1 vccd1 vccd1
+ _03712_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07303_ total_design.core.regFile.register\[23\]\[14\] net810 _02832_ _02833_ _02835_
+ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_117_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08283_ total_design.core.data_mem.last_read net998 vssd1 vssd1 vccd1 vccd1 _03675_
+ sky130_fd_sc_hd__nand2b_2
XFILLER_0_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout135_A _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload8 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_6
XFILLER_0_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07234_ _02755_ _02756_ _02769_ net683 total_design.core.regFile.register\[0\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__o32a_4
XFILLER_0_116_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08282__X _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11729__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09097__Y _04348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07165_ total_design.core.regFile.register\[1\]\[12\] net592 net570 total_design.core.regFile.register\[17\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__a22o_1
XANTENNA__10464__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1044_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07096_ _02637_ _02639_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06243__A _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1211_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout201 net204 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout212 _04721_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_1
Xfanout223 _04657_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout671_A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 net235 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_2
Xfanout245 net247 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout256 _04520_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout769_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09806_ net187 net2357 net439 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__mux2_1
Xfanout267 _04452_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout278 net279 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_2
Xfanout289 _04196_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_4
X_07998_ total_design.core.regFile.register\[30\]\[28\] net660 net603 total_design.core.regFile.register\[31\]\[28\]
+ _03490_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__a221o_1
XANTENNA__07581__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09737_ _04794_ _04957_ net320 vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06949_ total_design.core.regFile.register\[26\]\[8\] net645 net564 total_design.core.regFile.register\[3\]\[8\]
+ _02499_ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout936_A _05688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_66_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08125__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__A0 _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13125__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09668_ _04892_ _04893_ net704 vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07333__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08619_ total_design.lcd_display.cnt_20ms\[3\] _03910_ vssd1 vssd1 vccd1 vccd1 _03911_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06687__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10639__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ _04248_ _04272_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07521__B _03040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11630_ _05667_ net1690 net133 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06418__A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11561_ _05627_ net1663 net143 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13300_ clknet_leaf_142_clk _00767_ net1182 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10512_ net217 net2257 net480 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__mux2_1
X_14280_ net987 _01456_ net1084 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11492_ net1661 _05624_ net150 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13231_ clknet_leaf_147_clk _00698_ net1152 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10443_ net224 net2069 net383 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__mux2_1
XANTENNA__10374__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13162_ clknet_leaf_25_clk _00629_ net1106 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10374_ net237 net2364 net485 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__mux2_1
XANTENNA__06153__A total_design.core.ctrl.instruction\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12113_ net1525 net710 _05956_ _05969_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13093_ clknet_leaf_117_clk _00560_ net1161 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12145__B1 _05850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12044_ total_design.lcd_display.row_2\[82\] _05818_ _05846_ total_design.lcd_display.row_2\[98\]
+ _05903_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_72_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08364__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06299__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout790 net793 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_161_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12448__A1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13995_ clknet_leaf_89_clk _01175_ net1259 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_57_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_161_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08116__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12946_ clknet_leaf_145_clk _00413_ net1176 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07324__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06678__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10549__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12877_ clknet_leaf_0_clk _00344_ net1003 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11828_ total_design.lcd_display.cnt_20ms\[15\] total_design.lcd_display.cnt_20ms\[16\]
+ _05715_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__and3_1
XANTENNA__09365__A2_N _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14540__1312 vssd1 vssd1 vccd1 vccd1 net1312 _14540__1312/LO sky130_fd_sc_hd__conb_1
XANTENNA__06328__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14547_ total_design.lcd_display.lcd_en vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11759_ net97 net960 net293 total_design.core.data_bus_o\[31\] vssd1 vssd1 vccd1
+ vccd1 _01387_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09639__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14478_ clknet_leaf_38_clk _01545_ net1090 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10792__B total_design.core.data_bus_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload103 clknet_leaf_157_clk vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__bufinv_16
Xclkload114 clknet_leaf_164_clk vssd1 vssd1 vccd1 vccd1 clkload114/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_116_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload125 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 clkload125/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__10284__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13429_ clknet_leaf_158_clk _00896_ net1143 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06850__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload136 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 clkload136/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_116_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08262__B net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload147 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 clkload147/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_113_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload158 clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 clkload158/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_168_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload169 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 clkload169/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_168_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06602__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08970_ _04221_ _04222_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__nand2_1
XANTENNA__12136__B1 _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07921_ net749 _03421_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[26\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11409__A _05663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ total_design.core.regFile.register\[25\]\[25\] net648 net629 total_design.core.regFile.register\[5\]\[25\]
+ _03353_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__a221o_1
XANTENNA__06510__B net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09661__X _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06803_ total_design.core.regFile.register\[20\]\[5\] net672 net606 total_design.core.regFile.register\[15\]\[5\]
+ _02362_ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__a221o_1
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
X_07783_ total_design.core.regFile.register\[24\]\[24\] net791 _03285_ _03288_ vssd1
+ vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_48_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09522_ _04746_ _04754_ _04124_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__o21a_1
X_06734_ total_design.core.regFile.register\[28\]\[4\] net853 net758 total_design.core.regFile.register\[4\]\[4\]
+ _02297_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11111__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07622__A _03112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09453_ _03036_ net446 _04290_ _04664_ _04688_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__o221a_1
XANTENNA__06669__A2 _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10459__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06665_ total_design.core.regFile.register\[0\]\[2\] net682 _02226_ _02232_ vssd1
+ vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_148_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08404_ _03758_ _03759_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09384_ _04527_ _04622_ net329 vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__mux2_1
XANTENNA__06238__A net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06596_ total_design.core.regFile.register\[16\]\[1\] net744 net738 net736 vssd1
+ vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08335_ total_design.core.data_mem.data_write_adr_reg\[25\] net546 net538 total_design.core.data_mem.data_read_adr_reg\[25\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout517_A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout138_X net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08266_ net1396 net558 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[16\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_144_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07217_ total_design.core.regFile.register\[13\]\[13\] net666 net562 total_design.core.regFile.register\[3\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08197_ total_design.core.data_mem.data_write_adr_reg\[9\] total_design.core.data_mem.data_write_adr_reg\[8\]
+ total_design.core.data_mem.data_write_adr_reg\[11\] total_design.core.data_mem.data_write_adr_reg\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__or4_1
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08172__B _02893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09983__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07148_ _02666_ _02688_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_93_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07079_ total_design.core.regFile.register\[3\]\[10\] net865 net819 total_design.core.regFile.register\[17\]\[10\]
+ _02614_ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__a221o_1
XANTENNA__12127__B1 _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10090_ net269 net2643 net402 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__mux2_1
Xfanout1007 net1015 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06701__A _02266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1018 net1027 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__buf_2
Xfanout1029 net1036 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11350__A1 total_design.core.data_bus_o\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout841_X net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12800_ clknet_leaf_201_clk _00267_ net1003 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13780_ clknet_leaf_49_clk total_design.core.data_mem.stored_data_adr\[23\] net1103
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10992_ _05217_ _05221_ _05225_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__and3_1
X_12731_ clknet_leaf_145_clk _00198_ net1173 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10369__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12662_ clknet_leaf_153_clk _00129_ net1136 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06148__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14401_ clknet_leaf_45_clk _01538_ net1085 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11613_ _05645_ net1692 net137 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08806__B1 _02367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12593_ clknet_leaf_148_clk _00060_ net1148 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14332_ clknet_leaf_52_clk _01493_ net1093 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_137_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11544_ net1545 _05628_ net147 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07085__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08363__A _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14263_ clknet_leaf_101_clk _01442_ net1239 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.currentState\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09178__B _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11475_ net1595 _05636_ net154 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13214_ clknet_leaf_174_clk _00681_ net1053 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09893__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10426_ net163 net2408 net386 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14194_ clknet_leaf_79_clk _01374_ net1219 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13145_ clknet_leaf_197_clk _00612_ net1007 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10357_ net174 net2797 net489 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12118__B1 _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07793__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08810__B total_design.core.data_mem.data_cpu_i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ clknet_leaf_143_clk _00543_ net1175 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_163_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ net186 net2098 net498 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__mux2_1
X_12027_ total_design.lcd_display.row_1\[25\] _05838_ _05850_ total_design.lcd_display.row_2\[1\]
+ _05823_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__a221o_1
XANTENNA__06330__B _01905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06899__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09641__B net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13978_ clknet_leaf_84_clk _01158_ net1249 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09133__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12929_ clknet_leaf_164_clk _00396_ net1165 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10279__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08257__B net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_124_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06450_ total_design.core.ctrl.instruction\[20\] _02020_ _02021_ total_design.core.ctrl.instruction\[7\]
+ _02024_ vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[0\] sky130_fd_sc_hd__a221o_2
XFILLER_0_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06381_ total_design.core.regFile.register\[30\]\[0\] net927 net917 net947 vssd1
+ vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__and4_1
XFILLER_0_29_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08120_ total_design.core.regFile.register\[24\]\[31\] net791 net760 total_design.core.regFile.register\[21\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__a22o_1
XANTENNA__07076__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08051_ _03540_ _03542_ _03543_ _03545_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__or4_2
XFILLER_0_4_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06823__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06505__B net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07002_ total_design.core.regFile.register\[19\]\[9\] net642 net603 total_design.core.regFile.register\[31\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09222__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12109__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07784__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _02115_ _02187_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__nand2_1
XANTENNA__08328__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09525__A1 total_design.core.ctrl.instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07904_ total_design.core.regFile.register\[5\]\[26\] net629 net574 total_design.core.regFile.register\[24\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08884_ _04136_ _04137_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__nor2_1
XANTENNA__07536__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1007_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09391__X _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07835_ total_design.core.regFile.register\[24\]\[25\] net791 net760 total_design.core.regFile.register\[21\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__a22o_1
XANTENNA__07000__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11573__S net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__B _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07766_ total_design.core.regFile.register\[0\]\[23\] net682 _03266_ _03272_ vssd1
+ vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__o22a_4
XFILLER_0_79_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09505_ total_design.core.ctrl.instruction\[20\] net886 net754 total_design.core.data_cpu_o\[20\]
+ _04738_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a221o_1
X_06717_ total_design.core.regFile.register\[26\]\[3\] net646 _02281_ net687 vssd1
+ vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10189__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07697_ _03206_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[22\]
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout634_A _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09978__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09436_ _04277_ _04672_ _02337_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__o21ai_1
X_06648_ total_design.core.regFile.register\[2\]\[2\] net637 net621 total_design.core.regFile.register\[4\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09367_ _04601_ _04603_ _04606_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_23_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06579_ net903 _02019_ _01737_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08318_ net1463 net939 _03693_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[16\]
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_43_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07067__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12060__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ _04539_ _04540_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08249_ total_design.core.data_mem.state\[1\] _03657_ total_design.core.data_mem.state\[2\]
+ total_design.core.data_mem.state\[0\] vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__and4b_2
XFILLER_0_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06814__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09566__X _04797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ _05418_ _05508_ _05512_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__or3b_1
XFILLER_0_31_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10211_ _04720_ net2284 net391 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10652__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11191_ _05442_ _05446_ _05449_ _05439_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__09726__B _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10142_ net204 net2435 net400 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10073_ net209 net2173 net407 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__mux2_1
XANTENNA__07527__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12520__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ clknet_leaf_85_clk _01081_ net1249 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11483__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ clknet_leaf_60_clk _01040_ net1132 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07262__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13763_ clknet_leaf_60_clk total_design.core.data_mem.stored_data_adr\[6\] net1216
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10099__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10975_ _05233_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_139_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09888__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12714_ clknet_leaf_20_clk _00181_ net1050 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13694_ clknet_leaf_38_clk total_design.core.data_mem.stored_read_data\[1\] net1078
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12645_ clknet_leaf_119_clk _00112_ net1203 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07058__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12576_ clknet_leaf_194_clk _00043_ net1012 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14315_ clknet_leaf_63_clk _01476_ net1124 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_11527_ net1588 _05677_ net145 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__mux2_1
XANTENNA__06805__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold309 net66 vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14246_ clknet_leaf_109_clk _01426_ net1228 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11458_ net1622 _05635_ net155 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__mux2_1
XANTENNA__09204__B1 _04450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11658__S net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10409_ net233 net2197 net388 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__mux2_1
XANTENNA__10562__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14177_ clknet_leaf_112_clk net2705 net1208 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_2
X_11389_ _05578_ _05642_ _05647_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__o21a_2
X_13128_ clknet_leaf_24_clk _00595_ net1056 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07230__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13059_ clknet_leaf_15_clk _00526_ net1024 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1009 total_design.core.regFile.register\[13\]\[3\] vssd1 vssd1 vccd1 vccd1 net2325
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07620_ _03132_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_132_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07551_ total_design.core.regFile.register\[9\]\[19\] net851 net795 total_design.core.regFile.register\[11\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09798__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06502_ net746 net732 net726 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__and3_4
XFILLER_0_159_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07482_ total_design.core.regFile.register\[26\]\[18\] net644 net573 total_design.core.regFile.register\[24\]\[18\]
+ _03002_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07297__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09221_ _02537_ net504 net446 _02536_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__o22a_1
XFILLER_0_124_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12027__C1 _05823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06433_ total_design.core.regFile.register\[15\]\[0\] net846 _01983_ _01985_ _01991_
+ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_91_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09152_ total_design.core.data_cpu_o\[5\] net757 _04396_ _04400_ vssd1 vssd1 vccd1
+ vccd1 _04401_ sky130_fd_sc_hd__a211o_2
XANTENNA__09099__A _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07049__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12042__A2 _05839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06364_ net951 net950 total_design.core.ctrl.instruction\[20\] total_design.core.ctrl.instruction\[21\]
+ net952 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_161_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08103_ _03595_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__inv_2
XANTENNA__08797__A2 total_design.core.data_mem.data_cpu_i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_06295_ total_design.core.instr_mem.instruction_adr_i\[0\] total_design.core.instr_mem.instruction_adr_stored\[0\]
+ net984 vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__mux2_1
X_09083_ _02289_ net448 _04328_ _04333_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_141_Left_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08034_ _03526_ _03527_ _03528_ _03529_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold810 total_design.core.regFile.register\[2\]\[30\] vssd1 vssd1 vccd1 vccd1 net2126
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold821 total_design.core.regFile.register\[8\]\[0\] vssd1 vssd1 vccd1 vccd1 net2137
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11568__S net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold832 total_design.data_in_BUS\[22\] vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 total_design.core.regFile.register\[23\]\[27\] vssd1 vssd1 vccd1 vccd1 net2159
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_171_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10472__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold854 total_design.core.regFile.register\[8\]\[11\] vssd1 vssd1 vccd1 vccd1 net2170
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1124_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07757__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold865 total_design.core.regFile.register\[20\]\[29\] vssd1 vssd1 vccd1 vccd1 net2181
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 total_design.core.regFile.register\[27\]\[24\] vssd1 vssd1 vccd1 vccd1 net2192
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold887 total_design.core.regFile.register\[21\]\[21\] vssd1 vssd1 vccd1 vccd1 net2203
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold898 total_design.core.regFile.register\[7\]\[27\] vssd1 vssd1 vccd1 vccd1 net2214
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07221__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09985_ _04115_ _04982_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__nand2_4
XANTENNA_fanout584_A _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ _02117_ net505 net446 _02116_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__o22ai_1
XANTENNA__07509__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_186_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1510 total_design.core.regFile.register\[22\]\[3\] vssd1 vssd1 vccd1 vccd1 net2826
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1521 total_design.core.regFile.register\[10\]\[1\] vssd1 vssd1 vccd1 vccd1 net2837
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06401__D _01950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ _04120_ _04114_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__and2b_4
Xhold1532 total_design.core.regFile.register\[30\]\[15\] vssd1 vssd1 vccd1 vccd1 net2848
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout751_A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1543 total_design.core.regFile.register\[11\]\[7\] vssd1 vssd1 vccd1 vccd1 net2859
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_150_Left_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1554 total_design.data_in_BUS\[19\] vssd1 vssd1 vccd1 vccd1 net2870 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1565 total_design.data_in_BUS\[9\] vssd1 vssd1 vccd1 vccd1 net2881 sky130_fd_sc_hd__dlygate4sd3_1
X_07818_ _03303_ _03322_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_88_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08798_ _04034_ _04036_ _04042_ _04048_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__or4_1
XFILLER_0_93_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08609__C net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07749_ total_design.core.regFile.register\[19\]\[23\] net640 net620 total_design.core.regFile.register\[4\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__a22o_1
XANTENNA__10220__B net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10760_ _05020_ _01777_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07288__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12281__A2 _02893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09419_ _04122_ _04656_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10647__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10691_ _04991_ net532 vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__nand2_4
XANTENNA__09662__A_N _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_124_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12430_ _04113_ _04116_ _04972_ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_134_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12033__A2 _05834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06248__B1 _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12361_ _01622_ _01623_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14100_ clknet_leaf_98_clk _01280_ net1246 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07996__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11312_ _05569_ _05570_ net294 vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_160_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12292_ total_design.core.math.pc_val\[16\] net524 _06129_ _06130_ vssd1 vssd1 vccd1
+ vccd1 _01486_ sky130_fd_sc_hd__a22o_1
XANTENNA__07460__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_139_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11478__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14031_ clknet_leaf_83_clk _01211_ net1243 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_11243_ _05401_ _05499_ _05492_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_132_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10382__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11544__A1 _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07257__A _02770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ _05427_ _05429_ _05423_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06161__A total_design.core.ctrl.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_101_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10125_ net283 total_design.core.regFile.register\[18\]\[4\] net398 vssd1 vssd1 vccd1
+ vccd1 _00427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10056_ net277 net1953 net407 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__mux2_1
XANTENNA__11847__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06723__A1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13815_ clknet_leaf_72_clk total_design.core.data_mem.data_cpu_i\[24\] net1211 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10807__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07279__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13746_ clknet_leaf_113_clk total_design.core.data_mem.stored_write_data\[21\] net1207
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[21\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_174_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10958_ _05216_ _05188_ _05183_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__mux2_2
XFILLER_0_70_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08816__A _02263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13677_ clknet_leaf_49_clk total_design.core.data_mem.data_read_adr_i\[17\] net1101
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[17\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10557__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10889_ _05087_ _05123_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_14_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12628_ clknet_leaf_142_clk _00095_ net1175 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12024__A2 _05810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12559_ net1409 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11783__A1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold106 total_design.core.instr_mem.instruction_adr_stored\[20\] vssd1 vssd1 vccd1
+ vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07451__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold117 total_design.core.data_mem.data_bus_i_reg\[16\] vssd1 vssd1 vccd1 vccd1 net1433
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 total_design.core.instr_mem.instruction_adr_stored\[12\] vssd1 vssd1 vccd1
+ vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ clknet_leaf_48_clk _01409_ net1099 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dfrtp_1
Xhold139 total_design.core.data_mem.data_read_adr_reg2\[6\] vssd1 vssd1 vccd1 vccd1
+ net1455 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13062__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10292__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11535__A1 _05655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07739__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout608 net611 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_8
Xfanout619 _02068_ vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ net198 net2487 net444 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06982_ total_design.core.regFile.register\[31\]\[8\] net833 _02529_ _02532_ vssd1
+ vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__a211o_1
X_08721_ _03975_ _03980_ vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__nor2_1
Xfanout1190 net1200 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__clkbuf_2
X_08652_ total_design.lcd_display.cnt_500hz\[7\] _03936_ net712 vssd1 vssd1 vccd1
+ vccd1 _03937_ sky130_fd_sc_hd__a21boi_1
XANTENNA__07911__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07603_ total_design.core.regFile.register\[16\]\[20\] net854 net767 total_design.core.regFile.register\[7\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__a22o_1
X_08583_ _03769_ _03906_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[4\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07534_ total_design.core.regFile.register\[2\]\[19\] net637 net563 total_design.core.regFile.register\[3\]\[19\]
+ _03051_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__a221o_1
XANTENNA__12263__A2 _02796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10467__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07465_ net309 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[17\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1074_A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ _01754_ net753 _04450_ net904 _04447_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__o221a_2
XFILLER_0_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06416_ total_design.core.ctrl.instruction\[23\] net928 net919 net966 vssd1 vssd1
+ vccd1 vccd1 _01992_ sky130_fd_sc_hd__and4b_4
XFILLER_0_162_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12015__A2 _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07690__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07396_ total_design.core.regFile.register\[1\]\[16\] net828 net787 total_design.core.regFile.register\[13\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09135_ net328 _04267_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06347_ _01917_ _01920_ _01915_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07978__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09557__A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ _02240_ _04283_ _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_103_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06278_ total_design.core.data_adr_o\[3\] _01856_ net963 vssd1 vssd1 vccd1 vccd1
+ _01857_ sky130_fd_sc_hd__mux2_1
XANTENNA__07442__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08017_ total_design.core.regFile.register\[15\]\[29\] net846 net834 total_design.core.regFile.register\[10\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout799_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06650__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold640 total_design.core.regFile.register\[3\]\[26\] vssd1 vssd1 vccd1 vccd1 net1956
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08180__B _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11526__A1 _05626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold651 total_design.core.regFile.register\[10\]\[4\] vssd1 vssd1 vccd1 vccd1 net1967
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09991__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold662 total_design.core.regFile.register\[22\]\[5\] vssd1 vssd1 vccd1 vccd1 net1978
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold673 total_design.core.regFile.register\[20\]\[30\] vssd1 vssd1 vccd1 vccd1 net1989
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold684 total_design.core.regFile.register\[8\]\[29\] vssd1 vssd1 vccd1 vccd1 net2000
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold695 total_design.core.regFile.register\[30\]\[6\] vssd1 vssd1 vccd1 vccd1 net2011
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout587_X net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ net223 net2706 net420 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__mux2_1
X_08919_ net335 _03273_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__or2_1
X_09899_ net227 net2077 net428 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__mux2_1
Xhold1340 total_design.core.regFile.register\[29\]\[9\] vssd1 vssd1 vccd1 vccd1 net2656
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ total_design.keypad0.key_out\[10\] net529 net475 total_design.keypad0.key_out\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__a22o_1
Xhold1351 total_design.core.regFile.register\[0\]\[11\] vssd1 vssd1 vccd1 vccd1 net2667
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1362 total_design.core.regFile.register\[22\]\[27\] vssd1 vssd1 vccd1 vccd1 net2678
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1373 total_design.core.regFile.register\[19\]\[23\] vssd1 vssd1 vccd1 vccd1 net2689
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1384 total_design.core.regFile.register\[28\]\[4\] vssd1 vssd1 vccd1 vccd1 net2700
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07902__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1395 total_design.core.regFile.register\[30\]\[0\] vssd1 vssd1 vccd1 vccd1 net2711
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11861_ _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13600_ clknet_leaf_61_clk net1338 net1129 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _01728_ _05030_ net521 total_design.core.data_bus_o\[12\] _05028_ vssd1 vssd1
+ vccd1 vccd1 _05071_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11792_ net1767 net954 net301 _01804_ vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09655__B1 _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ clknet_leaf_143_clk _00998_ net1173 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10743_ net2879 net353 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10377__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13462_ clknet_leaf_152_clk _00929_ net1139 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12006__A2 _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07681__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06156__A total_design.core.ctrl.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10674_ net225 total_design.core.regFile.register\[2\]\[15\] net363 vssd1 vssd1 vccd1
+ vccd1 _00950_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12413_ net895 _01670_ net524 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13393_ clknet_leaf_151_clk _00860_ net1145 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12344_ net990 _01608_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07433__A2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12275_ total_design.core.math.pc_val\[15\] total_design.core.program_count.imm_val_reg\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11517__A1 _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14014_ clknet_leaf_101_clk _01194_ net1236 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[96\]
+ sky130_fd_sc_hd__dfrtp_1
X_11226_ _05484_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__inv_2
XANTENNA__08394__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ _05399_ _05406_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06944__A1 total_design.core.ctrl.instruction\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06944__B2 total_design.core.ctrl.instruction\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10108_ net204 net2147 net403 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__mux2_1
X_11088_ total_design.core.data_bus_o\[17\] net695 _05056_ _05299_ net517 vssd1 vssd1
+ vccd1 vccd1 _05347_ sky130_fd_sc_hd__a221o_1
X_10039_ net210 net2429 net411 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11671__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13729_ clknet_leaf_76_clk total_design.core.data_mem.stored_write_data\[4\] net1213
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10287__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07250_ total_design.core.regFile.register\[16\]\[13\] _01932_ net866 total_design.core.regFile.register\[3\]\[13\]
+ net694 vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06201_ total_design.core.data_adr_o\[29\] _01779_ net963 vssd1 vssd1 vccd1 vccd1
+ _01780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07181_ total_design.core.regFile.register\[3\]\[12\] net866 net854 total_design.core.regFile.register\[16\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11756__B2 total_design.core.data_bus_o\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09377__A _02818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06632__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11508__A1 _05636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09177__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout405 _04988_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_6
Xfanout416 _04983_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_6
X_09822_ net273 net2301 net437 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__mux2_1
Xfanout427 net429 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_8
Xfanout438 net441 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_6
XANTENNA__06935__A1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout449 net451 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_4
X_09753_ net257 net2111 net444 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__mux2_1
X_06965_ total_design.core.regFile.register\[3\]\[8\] net868 net817 total_design.core.regFile.register\[20\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout282_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08137__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ _00027_ _00026_ _03969_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__or3_1
XANTENNA__11147__A _05358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09684_ net507 _04909_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12484__A2 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06896_ total_design.core.regFile.register\[19\]\[7\] net640 net611 total_design.core.regFile.register\[18\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08635_ _03922_ _03923_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout547_A total_design.core.data_mem.next_write vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11581__S net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07360__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ total_design.data_in_BUS\[21\] net340 net719 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[21\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_81_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07517_ net308 _03035_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08497_ total_design.keypad0.key_out\[11\] _03848_ _03847_ vssd1 vssd1 vccd1 vccd1
+ _03849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08175__B _03040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout714_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09986__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07448_ total_design.core.regFile.register\[29\]\[17\] net798 net767 total_design.core.regFile.register\[7\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07663__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06407__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06871__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07379_ total_design.core.regFile.register\[23\]\[16\] net680 net672 total_design.core.regFile.register\[20\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout502_X net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11747__A1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ _02339_ net447 net289 _04366_ _04367_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__o221a_1
XANTENNA__07359__X total_design.core.data_mem.data_cpu_i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10390_ net173 net2199 net486 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__mux2_1
XANTENNA__06623__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09049_ _04178_ _04180_ net459 vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_4__f_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__06423__B net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12060_ total_design.lcd_display.row_2\[59\] net348 _05846_ total_design.lcd_display.row_2\[99\]
+ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a22o_1
Xhold470 _01364_ vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 total_design.lcd_display.row_2\[100\] vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout871_X net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold492 total_design.lcd_display.row_2\[79\] vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ _05248_ _05251_ _05253_ _05247_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__or4b_1
XANTENNA__08915__A2 _03322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10660__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout950 _01919_ vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_2
Xfanout961 _01770_ vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__buf_4
Xfanout972 total_design.core.ctrl.instruction\[6\] vssd1 vssd1 vccd1 vccd1 net972
+ sky130_fd_sc_hd__clkbuf_2
Xfanout983 net985 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_4
Xfanout994 net996 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ clknet_leaf_130_clk _00429_ net1199 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1170 total_design.core.regFile.register\[17\]\[16\] vssd1 vssd1 vccd1 vccd1 net2486
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ _05790_ total_design.data_from_keypad\[0\] net530 vssd1 vssd1 vccd1 vccd1
+ _01447_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11683__A0 _05651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1181 total_design.core.regFile.register\[1\]\[21\] vssd1 vssd1 vccd1 vccd1 net2497
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1192 total_design.core.regFile.register\[11\]\[26\] vssd1 vssd1 vccd1 vccd1 net2508
+ sky130_fd_sc_hd__dlygate4sd3_1
X_12893_ clknet_leaf_11_clk _00360_ net1025 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11491__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _05721_ _05730_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_16_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09628__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14563_ net35 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_1
X_11775_ net1693 net954 net301 _01836_ vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09896__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10726_ net2407 net354 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__and2_1
X_13514_ clknet_leaf_20_clk _00981_ net1050 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07654__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14494_ clknet_leaf_29_clk _01561_ net1073 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08851__A1 total_design.core.ctrl.instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_82_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06862__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13445_ clknet_leaf_116_clk _00912_ net1203 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10657_ net162 net2052 net477 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload15 clknet_leaf_200_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__inv_6
Xclkload26 clknet_leaf_179_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__bufinv_16
Xclkload37 clknet_leaf_191_clk vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__inv_8
X_13376_ clknet_leaf_3_clk _00843_ net1013 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07406__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10588_ net173 total_design.core.regFile.register\[5\]\[28\] net371 vssd1 vssd1 vccd1
+ vccd1 _00867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload48 clknet_leaf_172_clk vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__inv_6
XFILLER_0_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload59 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12327_ net899 _03138_ net522 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_77_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09159__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12258_ total_design.core.math.pc_val\[13\] total_design.core.program_count.imm_val_reg\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__and2_1
XANTENNA__11666__S net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ _05456_ _05463_ _05467_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__or3_1
XANTENNA__10570__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12189_ _06037_ _06038_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_166_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07445__A _02968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08119__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06750_ net721 _02312_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__nor2_1
XANTENNA__09867__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07327__D1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11674__A0 _05609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09660__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06681_ total_design.core.regFile.register\[25\]\[3\] net842 _02244_ _02247_ vssd1
+ vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08420_ total_design.keypad0.key_out\[5\] total_design.keypad0.key_out\[6\] total_design.keypad0.key_out\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__and3_1
XANTENNA__07893__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08351_ total_design.data_in_BUS\[0\] net512 _01904_ vssd1 vssd1 vccd1 vccd1 _03711_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_157_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07302_ total_design.core.regFile.register\[3\]\[14\] net866 net822 total_design.core.regFile.register\[17\]\[14\]
+ _02834_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__a221o_1
XANTENNA__06508__B net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08282_ total_design.core.data_mem.last_read net998 vssd1 vssd1 vccd1 vccd1 _03674_
+ sky130_fd_sc_hd__and2b_2
XFILLER_0_129_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload9 clknet_leaf_193_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__inv_6
X_07233_ total_design.core.regFile.register\[10\]\[13\] net616 _02763_ _02767_ _02768_
+ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06853__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11729__A1 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07179__X _02718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07164_ total_design.core.regFile.register\[5\]\[12\] net630 net587 total_design.core.regFile.register\[28\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07095_ _02587_ _02638_ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__or2_1
XANTENNA__08070__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1037_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11576__S net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 net204 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_1
XANTENNA_fanout497_A _05004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10480__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout213 net214 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout224 net227 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_2
Xfanout235 _04615_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1204_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout246 net247 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09805_ net191 net2756 net439 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__mux2_1
Xfanout257 net260 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07030__B1 _01995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout268 net271 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07997_ total_design.core.regFile.register\[26\]\[28\] net645 net638 total_design.core.regFile.register\[2\]\[28\]
+ _03493_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__a221o_1
Xfanout279 _04315_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_2
XANTENNA_fanout664_A net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06948_ total_design.core.regFile.register\[23\]\[8\] net680 net676 total_design.core.regFile.register\[22\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__a22o_1
X_09736_ _03644_ net505 net296 _04626_ _04958_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__o221a_1
Xclkbuf_4_12__f_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__11665__A0 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ _04871_ _04891_ _03509_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout831_A _01959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06879_ total_design.core.regFile.register\[17\]\[6\] net821 _02434_ _02435_ vssd1
+ vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout929_A net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08618_ total_design.lcd_display.cnt_20ms\[0\] total_design.lcd_display.cnt_20ms\[1\]
+ total_design.lcd_display.cnt_20ms\[2\] vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__and3_1
XANTENNA__12209__A2 _04450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ _03375_ net704 _04826_ net535 vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__a211o_1
XANTENNA__07884__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08549_ _03771_ _03800_ _03896_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12090__B1 _05912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11560_ _05677_ net1674 net141 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__mux2_1
XANTENNA__07636__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10511_ net214 net1934 net480 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06844__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11491_ net1612 _05635_ net151 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__mux2_1
XANTENNA__10655__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ clknet_leaf_189_clk _00697_ net1030 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442_ net234 net2688 net384 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09389__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13161_ clknet_leaf_178_clk _00628_ net1033 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10373_ net241 net2194 net485 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12112_ _05951_ _05965_ _05967_ _05968_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07817__X _03322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06721__X _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ clknet_leaf_108_clk _00559_ net1223 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11486__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12043_ total_design.lcd_display.row_1\[98\] _05810_ _05844_ total_design.lcd_display.row_2\[42\]
+ _05823_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__a221o_1
XANTENNA__10390__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07021__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout780 net782 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout791 net793 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_161_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13994_ clknet_leaf_86_clk _01174_ net1247 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11656__A0 _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ clknet_leaf_148_clk _00412_ net1146 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07875__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12876_ clknet_leaf_174_clk _00343_ net1054 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09746__A_N total_design.core.ctrl.instruction\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_158_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11827_ net1872 _05715_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06328__B net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12081__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11758_ net1864 net957 _05037_ _05695_ vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__a22o_1
X_14546_ total_design.lcd_display.lcd_rs vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07627__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10709_ net214 net2719 net357 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10565__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11689_ net2 net935 net878 net1852 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__o22a_1
X_14477_ clknet_leaf_40_clk _01544_ net1091 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09639__B _04866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10792__C total_design.core.data_bus_o\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload104 clknet_leaf_158_clk vssd1 vssd1 vccd1 vccd1 clkload104/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_144_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13428_ clknet_leaf_144_clk _00895_ net1176 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload115 clknet_leaf_165_clk vssd1 vssd1 vccd1 vccd1 clkload115/Y sky130_fd_sc_hd__inv_6
XFILLER_0_107_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload126 clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 clkload126/Y sky130_fd_sc_hd__inv_6
Xclkload137 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 clkload137/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_12_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload148 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 clkload148/Y sky130_fd_sc_hd__clkinv_8
Xclkload159 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 clkload159/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13359_ clknet_leaf_160_clk _00826_ net1150 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_max_cap348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08052__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07920_ _03418_ _03419_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__xnor2_4
XANTENNA__07012__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ total_design.core.regFile.register\[4\]\[25\] net621 net563 total_design.core.regFile.register\[3\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06510__C net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06802_ total_design.core.regFile.register\[11\]\[5\] net614 net587 total_design.core.regFile.register\[28\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__a22o_1
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_07782_ total_design.core.regFile.register\[2\]\[24\] net784 _03286_ _03287_ vssd1
+ vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__a211o_1
XANTENNA__11647__A0 _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09521_ net295 _04388_ _04753_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__o21ai_1
X_06733_ total_design.core.regFile.register\[18\]\[4\] net857 _01992_ total_design.core.regFile.register\[20\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09452_ net968 _03036_ _03037_ net537 vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__o211ai_1
X_06664_ _02214_ _02218_ _02228_ _02231_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__or4_1
XANTENNA__07866__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08403_ _03735_ _03738_ _03736_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_143_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09383_ _04572_ _04621_ net464 vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__mux2_1
X_06595_ total_design.core.regFile.register\[26\]\[1\] net746 net731 net723 vssd1
+ vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout245_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08334_ net1500 net938 _03701_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[24\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07079__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09389__X _04628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08815__A1 total_design.core.data_mem.data_cpu_i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08734__A _02395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08265_ net1504 net558 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[15\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__10475__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout412_A net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1154_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07216_ total_design.core.regFile.register\[16\]\[13\] net633 net628 total_design.core.regFile.register\[5\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06254__A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08196_ total_design.core.data_mem.data_write_adr_reg\[1\] total_design.core.data_mem.data_write_adr_reg\[0\]
+ total_design.core.data_mem.data_write_adr_reg\[3\] total_design.core.data_mem.data_write_adr_reg\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__or4_1
XFILLER_0_132_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07147_ net551 net300 _02646_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08043__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout200_X net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07251__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07078_ total_design.core.regFile.register\[1\]\[10\] net827 net775 total_design.core.regFile.register\[22\]\[10\]
+ _02622_ vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_93_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout781_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1008 net1015 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1019 net1021 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09543__A2 _04189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11638__A0 _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ _04600_ _04666_ _04935_ _04942_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__a211o_1
X_10991_ _05217_ _05224_ _05249_ _05222_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07306__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12730_ clknet_leaf_125_clk _00197_ net1189 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07857__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12661_ clknet_leaf_166_clk _00128_ net1157 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08793__A_N total_design.core.data_mem.data_cpu_i\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14400_ clknet_leaf_44_clk _01537_ net1085 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11612_ _05643_ net1719 net139 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__mux2_1
XANTENNA__09299__X _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12063__B1 _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12592_ clknet_leaf_182_clk _00059_ net1041 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08806__B2 _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14331_ clknet_leaf_39_clk _01492_ net1091 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11543_ net1666 _05612_ net145 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10385__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14262_ clknet_leaf_101_clk _01441_ net1239 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.currentState\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_11474_ net1657 _05652_ net155 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07490__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14134__RESET_B net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13213_ clknet_leaf_9_clk _00680_ net1019 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10425_ net165 net2149 net387 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14193_ clknet_leaf_80_clk _01373_ net1221 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13144_ clknet_leaf_136_clk _00611_ net1180 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07242__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06451__X _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10356_ net176 net2417 net489 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13075_ clknet_leaf_179_clk _00542_ net1035 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06170__Y _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10287_ net192 net2369 net498 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_163_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12026_ total_design.lcd_display.row_1\[113\] _05814_ _05852_ total_design.lcd_display.row_2\[9\]
+ _05886_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__a221o_1
XANTENNA__08742__B1 _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13977_ clknet_leaf_93_clk _01157_ net1253 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12928_ clknet_leaf_0_clk _00395_ net1003 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07848__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12859_ clknet_leaf_150_clk _00326_ net1147 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12054__B1 _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06380_ net926 net916 net946 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06808__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14529_ net1301 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_0_71_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08273__B net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08050_ total_design.core.regFile.register\[16\]\[29\] net632 net608 total_design.core.regFile.register\[18\]\[29\]
+ _03544_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__a221o_1
XANTENNA__07481__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07001_ _02547_ _02548_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08025__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09222__B2 _04466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08952_ _02115_ _02187_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__or2_1
XANTENNA__06521__B net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07903_ total_design.core.regFile.register\[25\]\[26\] net648 _03403_ net687 vssd1
+ vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__a211o_1
X_08883_ net334 _02666_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07834_ total_design.core.regFile.register\[23\]\[25\] net811 net795 total_design.core.regFile.register\[11\]\[25\]
+ _03337_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__a221o_1
X_07765_ _03268_ _03269_ _03270_ _03271_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout362_A net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06716_ total_design.core.regFile.register\[31\]\[3\] net602 net594 total_design.core.regFile.register\[8\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__a22o_1
X_09504_ net903 _04737_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07696_ total_design.core.regFile.register\[0\]\[22\] net875 _03191_ _03205_ vssd1
+ vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__o22ai_4
XANTENNA__07839__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09435_ net317 _04104_ _04484_ _04671_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__o31ai_1
X_06647_ total_design.core.regFile.register\[9\]\[2\] net664 net567 total_design.core.regFile.register\[12\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12045__B1 _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ _02841_ net508 net298 _04604_ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__o221a_1
X_06578_ total_design.core.ctrl.instruction\[3\] net906 vssd1 vssd1 vccd1 vccd1 _02150_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_23_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08317_ total_design.core.data_mem.data_write_adr_reg\[16\] net547 net539 total_design.core.data_mem.data_read_adr_reg\[16\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_43_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09297_ total_design.core.math.pc_val\[11\] _04516_ vssd1 vssd1 vccd1 vccd1 _04540_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09461__A1 total_design.core.ctrl.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08183__B _03421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09994__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08248_ net1428 net543 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[31\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_117_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06415__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08179_ net890 _03234_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[22\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10210_ net219 net2315 net389 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__mux2_1
X_11190_ _05442_ _05447_ _05440_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ net207 net2164 net399 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09516__A2 _03178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ net218 net2311 net406 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__mux2_1
X_13900_ clknet_leaf_73_clk _01080_ net1209 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[110\]
+ sky130_fd_sc_hd__dfrtp_1
X_13831_ clknet_leaf_78_clk _01039_ net1216 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07262__B _02796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13762_ clknet_leaf_61_clk total_design.core.data_mem.stored_data_adr\[5\] net1216
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[5\] sky130_fd_sc_hd__dfrtp_1
X_10974_ _05232_ _05195_ _05196_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_67_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12713_ clknet_leaf_3_clk _00180_ net1012 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13693_ clknet_leaf_40_clk total_design.core.data_mem.stored_read_data\[0\] net1092
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12036__B1 _05826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12644_ clknet_leaf_105_clk _00111_ net1233 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06446__X _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12575_ clknet_leaf_182_clk _00042_ net1043 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09452__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14314_ clknet_leaf_64_clk _01475_ net1124 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_11526_ net1519 _05626_ net147 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11457_ net1513 _05618_ net153 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__mux2_1
XANTENNA__08007__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14245_ clknet_leaf_104_clk _01425_ net1236 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09204__B2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10408_ net230 net1950 net388 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__mux2_1
X_14176_ clknet_leaf_114_clk _01356_ net1208 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfrtp_2
X_11388_ net304 net510 _05032_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__or3b_1
XFILLER_0_21_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10339_ net253 net2759 net488 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__mux2_1
X_13127_ clknet_leaf_176_clk _00594_ net1048 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06341__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13058_ clknet_leaf_127_clk _00525_ net1192 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11674__S net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12009_ _05864_ _05866_ _05868_ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_128_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06741__A2 _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07550_ total_design.core.regFile.register\[18\]\[19\] net858 net828 total_design.core.regFile.register\[1\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06501_ total_design.core.regFile.register\[15\]\[0\] net743 net733 net727 vssd1
+ vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__and4_1
XANTENNA__10825__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07481_ total_design.core.regFile.register\[29\]\[18\] net655 net569 total_design.core.regFile.register\[17\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09220_ net317 _04172_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06432_ total_design.core.regFile.register\[3\]\[0\] net865 _01962_ _01973_ _01939_
+ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__12027__B1 _05850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09151_ net905 _04399_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06363_ total_design.core.regFile.register\[26\]\[0\] net927 net917 net915 vssd1
+ vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__and4_1
XANTENNA__09443__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08102_ _03579_ _03580_ _03594_ net685 total_design.core.regFile.register\[0\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__o32a_4
XANTENNA__06516__B net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09082_ _04195_ _04332_ _04329_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07454__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06294_ net998 net997 total_design.core.data_adr_o\[0\] vssd1 vssd1 vccd1 vccd1 _01873_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08033_ total_design.core.regFile.register\[18\]\[29\] net857 net850 total_design.core.regFile.register\[9\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold800 total_design.core.regFile.register\[12\]\[5\] vssd1 vssd1 vccd1 vccd1 net2116
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 total_design.core.regFile.register\[7\]\[12\] vssd1 vssd1 vccd1 vccd1 net2127
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout208_A _04740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold822 total_design.core.regFile.register\[8\]\[22\] vssd1 vssd1 vccd1 vccd1 net2138
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 total_design.core.regFile.register\[10\]\[30\] vssd1 vssd1 vccd1 vccd1 net2149
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold844 total_design.core.regFile.register\[5\]\[25\] vssd1 vssd1 vccd1 vccd1 net2160
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 total_design.core.regFile.register\[27\]\[3\] vssd1 vssd1 vccd1 vccd1 net2171
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold866 total_design.core.regFile.register\[31\]\[26\] vssd1 vssd1 vccd1 vccd1 net2182
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08954__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold877 total_design.core.regFile.register\[5\]\[12\] vssd1 vssd1 vccd1 vccd1 net2193
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 total_design.core.regFile.register\[5\]\[26\] vssd1 vssd1 vccd1 vccd1 net2204
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 total_design.core.regFile.register\[6\]\[25\] vssd1 vssd1 vccd1 vccd1 net2215
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ _04112_ _04980_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout1117_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08935_ _01747_ _04123_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__or2_2
XANTENNA__11584__S net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1500 total_design.core.regFile.register\[25\]\[3\] vssd1 vssd1 vccd1 vccd1 net2816
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout577_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06980__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1511 total_design.core.regFile.register\[12\]\[8\] vssd1 vssd1 vccd1 vccd1 net2827
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 total_design.core.regFile.register\[18\]\[17\] vssd1 vssd1 vccd1 vccd1 net2838
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1533 total_design.core.regFile.register\[29\]\[8\] vssd1 vssd1 vccd1 vccd1 net2849
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08866_ _04118_ _04119_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__or2_1
XANTENNA__06717__C1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1544 total_design.core.regFile.register\[0\]\[30\] vssd1 vssd1 vccd1 vccd1 net2860
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1555 total_design.core.regFile.register\[28\]\[21\] vssd1 vssd1 vccd1 vccd1 net2871
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07817_ _03307_ _03308_ _03321_ net684 total_design.core.regFile.register\[0\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__o32a_4
Xhold1566 total_design.data_in_BUS\[24\] vssd1 vssd1 vccd1 vccd1 net2882 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_88_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08797_ _02565_ total_design.core.data_mem.data_cpu_i\[9\] _04044_ vssd1 vssd1 vccd1
+ vccd1 _04052_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_169_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08178__B _03187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06732__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09989__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ total_design.core.regFile.register\[31\]\[23\] net601 net593 total_design.core.regFile.register\[8\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07679_ total_design.core.regFile.register\[1\]\[22\] net828 net803 total_design.core.regFile.register\[8\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__a22o_1
XANTENNA__08906__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12018__B1 _05830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ _04655_ _04654_ _04650_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__nand3b_4
X_10690_ net162 net2424 net362 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_3__f_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09349_ net228 net2134 net453 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12360_ total_design.core.math.pc_val\[24\] net988 vssd1 vssd1 vccd1 vccd1 _01623_
+ sky130_fd_sc_hd__or2_1
X_11311_ _05564_ _05566_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12291_ net900 _02944_ net524 vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10663__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09198__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14030_ clknet_leaf_100_clk _01210_ net1229 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_11242_ _05401_ _05499_ _05492_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__or3b_1
XANTENNA__13708__RESET_B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12163__B total_design.core.data_access vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08945__B1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11173_ _05427_ _05429_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10124_ net269 net2023 net399 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__mux2_1
XANTENNA__11494__S net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06971__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10055_ net246 net1862 net409 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__mux2_1
XANTENNA__06723__A2 _02263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09899__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13814_ clknet_leaf_72_clk total_design.core.data_mem.data_cpu_i\[23\] net1205 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[23\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10807__A1 total_design.core.data_bus_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13745_ clknet_leaf_72_clk total_design.core.data_mem.stored_write_data\[20\] net1205
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[20\] sky130_fd_sc_hd__dfrtp_4
X_10957_ _05188_ _05190_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_123_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08816__B _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11480__A1 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07684__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13676_ clknet_leaf_56_clk total_design.core.data_mem.data_read_adr_i\[16\] net1113
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10888_ _05143_ _05144_ _05146_ _05127_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12627_ clknet_leaf_180_clk _00094_ net1041 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07436__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12558_ net1413 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11669__S net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11509_ net1619 _05609_ net151 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__mux2_1
XANTENNA__10573__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold107 total_design.core.math.pc_val\[26\] vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ net980 total_design.core.instr_mem.instruction_i\[8\] vssd1 vssd1 vccd1 vccd1
+ _01699_ sky130_fd_sc_hd__and2b_1
Xhold118 total_design.core.instr_mem.instruction_adr_stored\[30\] vssd1 vssd1 vccd1
+ vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold129 total_design.core.instr_mem.instruction_adr_stored\[17\] vssd1 vssd1 vccd1
+ vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14228_ clknet_leaf_48_clk _01408_ net1102 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08936__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14159_ clknet_leaf_31_clk _01339_ net1061 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout609 net611 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09663__A _04121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06981_ total_design.core.regFile.register\[14\]\[8\] net863 _02530_ _02531_ vssd1
+ vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_14__f_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06962__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ total_design.keypad0.counter\[0\] total_design.keypad0.counter\[1\] vssd1
+ vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12496__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1180 net1181 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__clkbuf_2
Xfanout1191 net1192 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__clkbuf_4
X_08651_ _03936_ net711 _03935_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__and3b_1
XANTENNA__06714__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ total_design.core.regFile.register\[24\]\[20\] net790 net783 total_design.core.regFile.register\[2\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__a22o_1
X_08582_ _03749_ net716 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[3\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_89_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07533_ total_design.core.regFile.register\[13\]\[19\] net667 net656 total_design.core.regFile.register\[29\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout158_A _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11471__A1 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07464_ total_design.core.regFile.register\[0\]\[17\] net873 _02980_ _02987_ vssd1
+ vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_48_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09203_ _04448_ _04449_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_85_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06415_ total_design.core.regFile.register\[22\]\[0\] net927 net917 net907 vssd1
+ vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__and4_1
XFILLER_0_91_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07395_ total_design.core.regFile.register\[6\]\[16\] net765 _02921_ vssd1 vssd1
+ vccd1 vccd1 _02922_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09134_ _04380_ _04381_ _04382_ net318 vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__o22a_1
X_06346_ _01914_ net950 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__nand2_1
XANTENNA__07427__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11774__A2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11579__S net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09065_ net333 net323 vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__nor2_1
X_06277_ total_design.core.instr_mem.instruction_adr_i\[3\] total_design.core.instr_mem.instruction_adr_stored\[3\]
+ net984 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10483__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08016_ net750 _03512_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[28\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 total_design.data_in_BUS\[18\] vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 total_design.core.regFile.register\[5\]\[7\] vssd1 vssd1 vccd1 vccd1 net1957
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08927__A0 _02917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold652 total_design.core.regFile.register\[7\]\[28\] vssd1 vssd1 vccd1 vccd1 net1968
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold663 total_design.core.regFile.register\[31\]\[5\] vssd1 vssd1 vccd1 vccd1 net1979
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold674 total_design.core.regFile.register\[16\]\[2\] vssd1 vssd1 vccd1 vccd1 net1990
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold685 total_design.core.regFile.register\[13\]\[5\] vssd1 vssd1 vccd1 vccd1 net2001
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 total_design.core.regFile.register\[28\]\[3\] vssd1 vssd1 vccd1 vccd1 net2012
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07645__X _03157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout861_A net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ net224 net2062 net420 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06953__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07364__Y _02893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ _04165_ _04171_ net325 vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__mux2_1
X_09898_ net234 net2807 net429 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__mux2_1
Xhold1330 total_design.core.regFile.register\[8\]\[31\] vssd1 vssd1 vccd1 vccd1 net2646
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1341 total_design.core.regFile.register\[16\]\[26\] vssd1 vssd1 vccd1 vccd1 net2657
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06201__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1352 total_design.core.regFile.register\[15\]\[8\] vssd1 vssd1 vccd1 vccd1 net2668
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1363 total_design.core.regFile.register\[21\]\[8\] vssd1 vssd1 vccd1 vccd1 net2679
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08849_ net968 net967 _04097_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__or3_4
XANTENNA__06705__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1374 total_design.core.data_bus_o\[0\] vssd1 vssd1 vccd1 vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1385 total_design.core.regFile.register\[2\]\[10\] vssd1 vssd1 vccd1 vccd1 net2701
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1396 total_design.core.regFile.register\[12\]\[29\] vssd1 vssd1 vccd1 vccd1 net2712
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11860_ total_design.lcd_display.currentState\[3\] _05724_ _05729_ _05744_ vssd1
+ vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_68_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10811_ net521 _05049_ _05064_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_0_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ net1812 net954 _05699_ _01838_ vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11462__A1 _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13530_ clknet_leaf_134_clk _00997_ net1190 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10742_ net2822 net353 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07130__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13461_ clknet_leaf_158_clk _00928_ net1143 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10673_ net232 net2571 net364 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_173_Right_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12412_ _04925_ _01669_ net993 vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13392_ clknet_leaf_184_clk _00859_ net1037 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11489__S net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12343_ _01595_ _01597_ _01598_ _01606_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__a211o_1
XANTENNA__10393__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12274_ total_design.core.math.pc_val\[15\] total_design.core.program_count.imm_val_reg\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11225_ _05362_ _05372_ _05378_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__and3_1
X_14013_ clknet_leaf_92_clk _01193_ net1259 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07197__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09483__A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ _05409_ _05410_ _05411_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10107_ net208 net2401 net405 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11087_ _05303_ net517 _05036_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__or3b_1
XANTENNA__12478__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10038_ net216 net2709 net410 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_170_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10568__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ _05746_ _05749_ _05798_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__or3_4
XFILLER_0_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11453__A1 _05630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13728_ clknet_leaf_76_clk total_design.core.data_mem.stored_write_data\[3\] net1214
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07657__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07121__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13659_ clknet_leaf_54_clk total_design.core.data_mem.data_write_adr_i\[31\] net1113
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[31\] sky130_fd_sc_hd__dfrtp_1
X_06200_ total_design.core.instr_mem.instruction_adr_i\[29\] total_design.core.instr_mem.instruction_adr_stored\[29\]
+ net983 vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_185_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07180_ total_design.core.regFile.register\[17\]\[12\] net822 net785 total_design.core.regFile.register\[2\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11756__A2 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07188__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout406 net409 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_8
X_09821_ net259 net2139 net437 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__mux2_1
Xfanout417 _04983_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_4
Xfanout428 net429 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_8
Xfanout439 net441 vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_6
XANTENNA__06935__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ net280 net2490 net442 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_123_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06964_ _02500_ _02501_ _02514_ net685 total_design.core.regFile.register\[0\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__o32a_4
XTAP_TAPCELL_ROW_33_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08703_ _00025_ _00024_ _00023_ _03968_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__or4_1
X_06895_ _02399_ _02440_ _02439_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__a21bo_2
X_09683_ _01757_ net753 _02897_ _04904_ _04908_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__o2111ai_4
XANTENNA__11862__S net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06699__A1 total_design.core.ctrl.instruction\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07896__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06699__B2 total_design.core.ctrl.instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08634_ total_design.lcd_display.cnt_500hz\[7\] total_design.lcd_display.cnt_500hz\[6\]
+ total_design.lcd_display.cnt_500hz\[9\] total_design.lcd_display.cnt_500hz\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__or4_1
XFILLER_0_90_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08737__A _02796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07360__A2 total_design.core.data_mem.data_cpu_i\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_138_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09637__A1 total_design.core.ctrl.instruction\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10478__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ total_design.data_in_BUS\[20\] net341 net719 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[20\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_138_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09637__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout442_A _04969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11444__A1 _05612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07516_ net308 _03035_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__or2_1
X_08496_ total_design.keypad0.key_out\[11\] _03808_ vssd1 vssd1 vccd1 vccd1 _03848_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07112__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11995__A2 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07447_ total_design.core.regFile.register\[19\]\[17\] net823 net802 total_design.core.regFile.register\[8\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_170_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_170_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_80_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout707_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07378_ total_design.core.regFile.register\[25\]\[16\] net649 net609 total_design.core.regFile.register\[18\]\[16\]
+ _02899_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_3_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11747__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06329_ net997 _01906_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__nor2_1
X_09117_ net969 _02339_ _02340_ _04100_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_115_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08073__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07088__A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09048_ _04299_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06423__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold460 total_design.lcd_display.row_2\[43\] vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold471 net58 vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 net70 vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08376__A1 _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11010_ _05248_ _05251_ _05254_ _05256_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_129_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07179__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold493 net65 vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09507__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout864_X net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 _03675_ vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06926__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout951 _01916_ vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__buf_2
Xfanout962 _01770_ vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout973 total_design.core.ctrl.instruction\[5\] vssd1 vssd1 vccd1 vccd1 net973
+ sky130_fd_sc_hd__buf_4
Xfanout984 net985 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__buf_4
Xfanout995 net996 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ clknet_leaf_121_clk _00428_ net1170 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1160 total_design.core.ctrl.instruction\[1\] vssd1 vssd1 vccd1 vccd1 net2476
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 total_design.core.regFile.register\[29\]\[22\] vssd1 vssd1 vccd1 vccd1 net2487
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ _03908_ _05776_ _05779_ _05788_ _05789_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__a311o_1
Xhold1182 total_design.core.regFile.register\[17\]\[8\] vssd1 vssd1 vccd1 vccd1 net2498
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07887__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 total_design.core.regFile.register\[17\]\[2\] vssd1 vssd1 vccd1 vccd1 net2509
+ sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ clknet_leaf_31_clk _00359_ net1060 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07351__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _05728_ _05729_ _05727_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__o21a_1
XANTENNA__10388__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08366__B net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11435__A1 _05655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07639__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14562_ net1282 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
X_11774_ net1795 net955 net301 _01849_ vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13513_ clknet_leaf_178_clk _00980_ net1047 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10725_ total_design.core.regFile.register\[0\]\[0\] net354 vssd1 vssd1 vccd1 vccd1
+ _00999_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_161_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_161_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14493_ clknet_leaf_27_clk _01560_ net1077 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07154__A_N total_design.core.ctrl.instruction\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08851__A2 total_design.core.ctrl.instruction\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_126_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13444_ clknet_leaf_107_clk _00911_ net1223 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10656_ net165 net2445 net478 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11520__B _05478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload16 clknet_leaf_201_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__clkinvlp_4
X_13375_ clknet_leaf_181_clk _00842_ net1043 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload27 clknet_leaf_180_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__bufinv_16
X_10587_ net179 net2046 net372 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__mux2_1
XANTENNA__06173__Y _01755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload38 clknet_leaf_192_clk vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_118_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload49 clknet_leaf_173_clk vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__inv_6
XANTENNA__06614__B _02182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12326_ net990 _01590_ _01591_ _01592_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a31o_1
XANTENNA__07811__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12257_ total_design.core.math.pc_val\[13\] total_design.core.program_count.imm_val_reg\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07285__X _02818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09564__B1 _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ _05455_ _05465_ _05450_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_142_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12188_ total_design.core.math.pc_val\[5\] total_design.core.program_count.imm_val_reg\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_166_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06917__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11139_ _05395_ _05397_ _05391_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07590__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12605__RESET_B net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11682__S net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06680_ total_design.core.regFile.register\[15\]\[3\] net847 _02245_ _02246_ vssd1
+ vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__a211o_1
XANTENNA__07342__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10298__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08350_ total_design.core.mem_ctrl.next_next_data_read _01774_ vssd1 vssd1 vccd1
+ vccd1 _03710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11426__A1 _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07301_ total_design.core.regFile.register\[15\]\[14\] net849 net841 total_design.core.regFile.register\[30\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06508__C net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08281_ net1369 net557 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[31\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__06302__B1 _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_152_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_152_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07232_ total_design.core.regFile.register\[18\]\[13\] net611 net588 total_design.core.regFile.register\[28\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13464__RESET_B net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11729__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07163_ total_design.core.regFile.register\[11\]\[12\] net612 net577 total_design.core.regFile.register\[27\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07094_ _02496_ _02539_ _02585_ _02536_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__o211a_1
XANTENNA__07802__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11857__S net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_2
Xfanout214 net215 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06540__A _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout392_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout225 net227 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_2
Xfanout236 net239 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_2
X_09804_ net195 net2636 net438 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__mux2_1
Xfanout247 _04281_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_31_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout258 net260 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_2
Xfanout269 net271 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_2
X_07996_ total_design.core.regFile.register\[11\]\[28\] net613 net568 total_design.core.regFile.register\[12\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__a22o_1
XANTENNA__07581__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09735_ net305 _03643_ net448 vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__or3_1
X_06947_ total_design.core.regFile.register\[13\]\[8\] net668 net638 total_design.core.regFile.register\[2\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11592__S net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout657_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09666_ _04871_ _04891_ _03509_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__o21bai_2
X_06878_ total_design.core.regFile.register\[31\]\[6\] net833 net825 total_design.core.regFile.register\[19\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07333__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08617_ total_design.lcd_display.cnt_20ms\[0\] total_design.lcd_display.cnt_20ms\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09597_ _04824_ _04825_ net707 vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout824_A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08186__B _03559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09997__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07090__B _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10001__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ total_design.keypad0.key_out\[13\] net932 net931 vssd1 vssd1 vccd1 vccd1
+ _03896_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08479_ _03830_ _03831_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_143_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_143_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08914__B _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10510_ net223 net2584 net482 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11490_ net1554 _05618_ net149 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10441_ net228 net1896 net381 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08046__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09243__C1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10372_ net255 net2226 net484 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13160_ clknet_leaf_170_clk _00627_ net1159 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout981_X net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12111_ total_design.lcd_display.row_2\[101\] _05846_ _05912_ vssd1 vssd1 vccd1 vccd1
+ _05968_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13091_ clknet_leaf_5_clk _00558_ net1022 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10671__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12145__A2 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ total_design.lcd_display.row_1\[58\] _05839_ _05849_ total_design.lcd_display.row_2\[50\]
+ _05901_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__a221o_1
Xhold290 total_design.lcd_display.row_1\[78\] vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout770 _01996_ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__buf_4
Xfanout781 net782 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_4
Xfanout792 net793 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__buf_4
X_13993_ clknet_leaf_94_clk _01173_ net1255 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_161_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ clknet_leaf_182_clk _00411_ net1041 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07324__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12875_ clknet_leaf_115_clk _00342_ net1202 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11826_ _05715_ net1880 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__nor2_1
XANTENNA__06328__C _01905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14545_ net1267 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_134_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_134_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11757_ net94 net960 net293 total_design.core.data_bus_o\[29\] vssd1 vssd1 vccd1
+ vccd1 _01385_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10708_ net221 net2534 net359 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14476_ clknet_leaf_40_clk _01543_ net1090 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_11688_ total_design.bus_full net937 wishbone.prev_BUSY_O vssd1 vssd1 vccd1 vccd1
+ _05691_ sky130_fd_sc_hd__or3b_1
XFILLER_0_71_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13427_ clknet_leaf_190_clk _00894_ net1034 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload105 clknet_leaf_159_clk vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__clkinv_8
Xclkload116 clknet_leaf_166_clk vssd1 vssd1 vccd1 vccd1 clkload116/Y sky130_fd_sc_hd__clkinv_2
X_10639_ net230 net1981 net476 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload127 clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 clkload127/Y sky130_fd_sc_hd__inv_6
XFILLER_0_141_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09785__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06344__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload138 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 clkload138/Y sky130_fd_sc_hd__clkinv_4
Xclkload149 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 clkload149/Y sky130_fd_sc_hd__inv_6
X_13358_ clknet_leaf_186_clk _00825_ net1030 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11592__A0 _05626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11677__S net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12309_ net992 _04696_ _01577_ net894 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__o211a_1
XANTENNA__10581__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13289_ clknet_leaf_16_clk _00756_ net1023 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12136__A2 _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07850_ total_design.core.regFile.register\[9\]\[25\] net664 net571 total_design.core.regFile.register\[17\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__a22o_1
XANTENNA__11409__C _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07563__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06801_ total_design.core.regFile.register\[6\]\[5\] net584 net575 total_design.core.regFile.register\[24\]\[5\]
+ _02360_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__a221o_1
XANTENNA__06510__D net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07781_ total_design.core.regFile.register\[3\]\[24\] net867 net847 total_design.core.regFile.register\[15\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_09520_ _04196_ _04751_ _04752_ _04748_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__o211a_1
X_06732_ total_design.core.regFile.register\[3\]\[4\] net865 net854 total_design.core.regFile.register\[16\]\[4\]
+ _02295_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a221o_1
X_09451_ net312 _04193_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__nand2_2
X_06663_ _02216_ _02217_ _02229_ _02230_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06519__B _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08402_ total_design.keypad0.key_out\[10\] _03757_ vssd1 vssd1 vccd1 vccd1 _03758_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06594_ total_design.core.regFile.register\[5\]\[1\] net741 net734 net728 vssd1 vssd1
+ vccd1 vccd1 _02165_ sky130_fd_sc_hd__and4_1
X_09382_ _04219_ _04222_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ total_design.core.data_mem.data_write_adr_reg\[24\] net546 net538 total_design.core.data_mem.data_read_adr_reg\[24\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_125_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout140_A _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08815__A2 _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08734__B _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout238_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08264_ net1354 net559 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[14\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__06535__A total_design.core.data_mem.data_cpu_i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07215_ _02742_ _02745_ _02740_ vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_15_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08028__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08195_ total_design.core.data_mem.data_write_adr_reg\[5\] total_design.core.data_mem.data_write_adr_reg\[4\]
+ total_design.core.data_mem.data_write_adr_reg\[7\] total_design.core.data_mem.data_write_adr_reg\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__or4_1
XFILLER_0_85_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07146_ net551 net300 _02646_ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__o21a_1
XANTENNA__11583__A0 _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11587__S net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07077_ total_design.core.regFile.register\[31\]\[10\] net831 _01980_ total_design.core.regFile.register\[12\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__a22o_1
XANTENNA__10491__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12127__A2 _05830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1009 net1015 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout774_A _01994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07554__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout941_A _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06762__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ total_design.core.regFile.register\[10\]\[28\] net835 net781 total_design.core.regFile.register\[27\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08909__B _03595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09718_ _04195_ _04936_ _04938_ _04941_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10990_ _05217_ _05225_ _05221_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__a21o_1
XANTENNA__07306__A2 total_design.core.data_mem.data_cpu_i\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09649_ _04875_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout827_X net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ clknet_leaf_140_clk _00127_ net1182 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11611_ _05648_ net1724 net137 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10666__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12591_ clknet_leaf_146_clk _00058_ net1153 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_116_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14330_ clknet_leaf_39_clk _01491_ net1091 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_11542_ net1557 _05609_ net147 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08019__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14261_ clknet_leaf_102_clk _01440_ net1239 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.currentState\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_11473_ net1544 _05613_ net153 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13212_ clknet_leaf_10_clk _00679_ net1021 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10424_ net171 net2073 net385 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__mux2_1
X_14192_ clknet_leaf_80_clk _01372_ net1221 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11574__A0 _05636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11497__S net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ clknet_leaf_166_clk _00610_ net1157 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10355_ net182 net2081 net489 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12118__A2 _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07793__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13074_ clknet_leaf_137_clk _00541_ net1179 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10286_ net195 net1926 net496 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12025_ total_design.lcd_display.row_2\[25\] _05832_ _05844_ total_design.lcd_display.row_2\[41\]
+ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a22o_1
XANTENNA__08742__A1 _03559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09491__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13976_ clknet_leaf_109_clk _01156_ net1225 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12927_ clknet_leaf_182_clk _00394_ net1043 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12858_ clknet_leaf_132_clk _00325_ net1196 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11809_ net1816 _05705_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10576__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_107_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12789_ clknet_leaf_158_clk _00256_ net1155 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_1_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14528_ net1300 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_0_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14459_ clknet_leaf_39_clk net1408 net1095 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09207__C1 _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07000_ total_design.core.regFile.register\[13\]\[9\] net668 net638 total_design.core.regFile.register\[2\]\[9\]
+ _02545_ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__a221o_1
XANTENNA__12357__A2 _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06505__D net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11565__A0 _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09222__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12109__A2 _05810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07784__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08951_ _01922_ _02445_ _04202_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__or3_4
XANTENNA__06521__C net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07902_ total_design.core.regFile.register\[8\]\[26\] net594 net563 total_design.core.regFile.register\[3\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__a22o_1
X_08882_ net470 _02613_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__nor2_1
XANTENNA__07536__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ total_design.core.regFile.register\[26\]\[25\] net870 net784 total_design.core.regFile.register\[2\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__a22o_1
XANTENNA__06744__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07764_ total_design.core.regFile.register\[30\]\[23\] net659 net608 total_design.core.regFile.register\[18\]\[23\]
+ _03257_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09503_ _04735_ _04736_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__or2_1
X_06715_ _02273_ _02275_ _02277_ _02279_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__or4_1
XFILLER_0_154_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07695_ total_design.core.regFile.register\[21\]\[22\] net760 _03192_ _03195_ _03204_
+ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout355_A _05018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07920__Y _03421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ net312 _04104_ _04670_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06646_ total_design.core.regFile.register\[25\]\[2\] net648 net602 total_design.core.regFile.register\[31\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10486__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09365_ _02839_ _04188_ net504 _02840_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout143_X net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06577_ _01735_ net903 vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__nor2_4
XFILLER_0_75_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1264_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08316_ net1456 net940 _03692_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[15\]
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_23_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09296_ total_design.core.math.pc_val\[11\] _04516_ vssd1 vssd1 vccd1 vccd1 _04539_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_43_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08247_ net1495 net542 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[30\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_145_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06415__D net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ net890 _03187_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[21\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11556__A0 _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout891_A _02022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07129_ total_design.core.regFile.register\[29\]\[11\] net801 _02667_ _02670_ vssd1
+ vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10140_ net209 net2553 net400 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__mux2_1
XANTENNA__06204__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ net214 net2747 net406 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__mux2_1
XANTENNA__07527__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_X net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06735__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13830_ clknet_leaf_77_clk _01038_ net1216 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13761_ clknet_leaf_61_clk total_design.core.data_mem.stored_data_adr\[4\] net1216
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[4\] sky130_fd_sc_hd__dfrtp_1
X_10973_ _05180_ _05195_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12712_ clknet_leaf_170_clk _00179_ net1159 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ clknet_leaf_47_clk net998 net1098 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.last_read
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12643_ clknet_leaf_5_clk _00110_ net1022 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10396__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ clknet_leaf_175_clk _00041_ net1053 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14313_ clknet_leaf_64_clk _01474_ net1124 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11525_ net1761 _05624_ net146 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09486__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14244_ clknet_leaf_104_clk _01424_ net1236 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11456_ net1702 _05621_ net155 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__mux2_1
XANTENNA__09204__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_944 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10407_ net236 net2565 net388 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__mux2_1
X_14175_ clknet_leaf_48_clk _01355_ net1099 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfrtp_2
XANTENNA__07718__B _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11387_ _05033_ _05610_ _05642_ _05587_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__o22a_4
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06622__B net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07766__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13126_ clknet_leaf_199_clk _00593_ net1001 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10338_ net251 net2737 net490 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__mux2_1
XANTENNA__06974__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13057_ clknet_leaf_121_clk _00524_ net1170 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10269_ net272 net1899 net499 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12008_ _05801_ _05824_ _05859_ _05869_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__or4_1
XFILLER_0_108_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13959_ clknet_leaf_82_clk _01139_ net1220 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06500_ net741 net733 net726 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__and3_1
X_07480_ total_design.core.regFile.register\[25\]\[18\] net647 net628 total_design.core.regFile.register\[5\]\[18\]
+ _02997_ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06431_ total_design.core.regFile.register\[28\]\[0\] net853 _01971_ _01977_ _01989_
+ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_9_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06356__Y _01932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09150_ _04397_ _04398_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06362_ net925 net917 net914 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__and3_1
XFILLER_0_161_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08101_ total_design.core.regFile.register\[31\]\[30\] net603 _03587_ _03592_ _03593_
+ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06516__C net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06293_ _01870_ _01855_ _01858_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__or3b_2
X_09081_ net323 _04331_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08032_ total_design.core.regFile.register\[16\]\[29\] _01932_ net775 total_design.core.regFile.register\[22\]\[29\]
+ net691 vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold801 total_design.core.regFile.register\[4\]\[0\] vssd1 vssd1 vccd1 vccd1 net2117
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold812 total_design.core.regFile.register\[25\]\[25\] vssd1 vssd1 vccd1 vccd1 net2128
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold823 total_design.core.regFile.register\[27\]\[5\] vssd1 vssd1 vccd1 vccd1 net2139
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold834 total_design.core.regFile.register\[15\]\[6\] vssd1 vssd1 vccd1 vccd1 net2150
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 total_design.core.regFile.register\[24\]\[20\] vssd1 vssd1 vccd1 vccd1 net2161
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07757__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold856 total_design.core.regFile.register\[5\]\[15\] vssd1 vssd1 vccd1 vccd1 net2172
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold867 total_design.core.regFile.register\[20\]\[4\] vssd1 vssd1 vccd1 vccd1 net2183
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 total_design.core.regFile.register\[11\]\[11\] vssd1 vssd1 vccd1 vccd1 net2194
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ net161 net2810 net419 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__mux2_1
Xhold889 total_design.core.regFile.register\[30\]\[17\] vssd1 vssd1 vccd1 vccd1 net2205
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06965__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10761__B2 total_design.core.data_access vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08934_ _01747_ _04123_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__nor2_2
XFILLER_0_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07509__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1501 total_design.core.regFile.register\[11\]\[29\] vssd1 vssd1 vccd1 vccd1 net2817
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12502__A2 total_design.core.ctrl.instruction\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1512 total_design.core.regFile.register\[20\]\[12\] vssd1 vssd1 vccd1 vccd1 net2828
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08865_ total_design.core.ctrl.instruction\[9\] total_design.core.ctrl.instruction\[10\]
+ net556 vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__o21a_1
Xhold1523 total_design.data_in_BUS\[21\] vssd1 vssd1 vccd1 vccd1 net2839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 total_design.core.regFile.register\[12\]\[15\] vssd1 vssd1 vccd1 vccd1 net2850
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11166__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1545 total_design.core.regFile.register\[17\]\[5\] vssd1 vssd1 vccd1 vccd1 net2861
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07816_ total_design.core.regFile.register\[29\]\[24\] net656 _03314_ _03319_ _03320_
+ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__a2111o_1
Xhold1556 total_design.core.regFile.register\[22\]\[28\] vssd1 vssd1 vccd1 vccd1 net2872
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1567 total_design.lcd_display.row_2\[34\] vssd1 vssd1 vccd1 vccd1 net2883 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_88_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08796_ _04047_ _04050_ _04049_ _04035_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_88_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07747_ _03183_ _03230_ _03232_ _03227_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07678_ total_design.core.regFile.register\[18\]\[22\] net858 net784 total_design.core.regFile.register\[2\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09417_ total_design.core.ctrl.instruction\[16\] net886 net754 total_design.core.data_cpu_o\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__a22o_1
X_06629_ total_design.core.regFile.register\[3\]\[2\] net867 net846 total_design.core.regFile.register\[15\]\[2\]
+ _02198_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout904_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09348_ net506 _04588_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_134_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09279_ _04500_ _04521_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08922__B _03112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11310_ _05531_ _05568_ _05562_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07996__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12290_ net993 _06126_ _06127_ _06128_ vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_151_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11241_ _05400_ _05499_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09198__B2 _04443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07748__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11172_ _05427_ _05430_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__and2_1
XANTENNA__06956__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ net278 net2251 net398 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__mux2_1
XANTENNA__07825__Y _03330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ net285 total_design.core.regFile.register\[20\]\[0\] net409 vssd1 vssd1 vccd1
+ vccd1 _00359_ sky130_fd_sc_hd__mux2_1
XANTENNA__06708__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11701__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06217__D_N _01795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07381__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13813_ clknet_leaf_111_clk total_design.core.data_mem.data_cpu_i\[22\] net1207 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[22\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13744_ clknet_leaf_112_clk total_design.core.data_mem.stored_write_data\[19\] net1207
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[19\] sky130_fd_sc_hd__dfrtp_1
X_10956_ _05213_ _05214_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06457__X _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07133__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13675_ clknet_leaf_58_clk total_design.core.data_mem.data_read_adr_i\[15\] net1118
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[15\] sky130_fd_sc_hd__dfrtp_1
X_10887_ _05121_ _05125_ _05087_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_155_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12626_ clknet_leaf_145_clk _00093_ net1179 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11768__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12180__C_N net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12557_ net1445 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_171_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10440__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ net1642 _05636_ net150 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_91_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12488_ net979 total_design.core.ctrl.instruction\[7\] net883 _01698_ vssd1 vssd1
+ vccd1 vccd1 _01546_ sky130_fd_sc_hd__a22o_1
Xhold108 total_design.core.instr_mem.instruction_adr_stored\[29\] vssd1 vssd1 vccd1
+ vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ clknet_leaf_49_clk _01407_ net1103 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__dfrtp_1
Xhold119 total_design.core.data_mem.data_read_adr_reg2\[21\] vssd1 vssd1 vccd1 vccd1
+ net1435 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ net1548 _05657_ net159 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07739__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14158_ clknet_leaf_31_clk _01338_ net1061 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06947__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13109_ clknet_leaf_160_clk _00576_ net1150 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09663__B _04889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14089_ clknet_leaf_93_clk _01269_ net1255 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_06980_ total_design.core.regFile.register\[10\]\[8\] net835 net769 total_design.core.regFile.register\[7\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1170 net1171 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__clkbuf_4
Xfanout1181 net1201 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__buf_2
X_08650_ total_design.lcd_display.cnt_500hz\[5\] total_design.lcd_display.cnt_500hz\[6\]
+ _03931_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__and3_1
Xfanout1192 net1194 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11417__C _05478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07372__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07601_ total_design.core.regFile.register\[30\]\[20\] net838 net834 total_design.core.regFile.register\[10\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__a22o_1
XANTENNA__07911__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08581_ _03734_ _03906_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[2\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07532_ _03048_ _03049_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07470__Y _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07463_ _02981_ _02983_ _02984_ _02986_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ total_design.core.math.pc_val\[5\] total_design.core.math.pc_val\[6\] _04371_
+ total_design.core.math.pc_val\[7\] vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09678__X _04904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06414_ net928 net917 net907 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__and3_4
XFILLER_0_85_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07394_ total_design.core.regFile.register\[25\]\[16\] net843 net825 total_design.core.regFile.register\[19\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_40_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11759__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ _04224_ _04259_ net323 vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__mux2_1
X_06345_ net971 net952 total_design.core.ctrl.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ _01921_ sky130_fd_sc_hd__and3b_1
XFILLER_0_161_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07978__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06276_ _01854_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__inv_2
X_09064_ net276 net1910 net453 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06543__A _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08015_ _03510_ _03511_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__or2_4
XFILLER_0_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06650__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold620 total_design.core.regFile.register\[31\]\[6\] vssd1 vssd1 vccd1 vccd1 net1936
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 total_design.core.regFile.register\[19\]\[7\] vssd1 vssd1 vccd1 vccd1 net1947
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold642 total_design.core.regFile.register\[27\]\[26\] vssd1 vssd1 vccd1 vccd1 net1958
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08927__A1 _02968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold653 total_design.core.regFile.register\[21\]\[0\] vssd1 vssd1 vccd1 vccd1 net1969
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 total_design.core.regFile.register\[29\]\[25\] vssd1 vssd1 vccd1 vccd1 net1980
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold675 total_design.core.regFile.register\[10\]\[17\] vssd1 vssd1 vccd1 vccd1 net1991
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold686 total_design.core.regFile.register\[18\]\[0\] vssd1 vssd1 vccd1 vccd1 net2002
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11595__S net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout687_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold697 total_design.core.regFile.register\[24\]\[9\] vssd1 vssd1 vccd1 vccd1 net2013
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ net232 net1961 net421 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1015_X net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ _04170_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__inv_2
X_09897_ net228 net1907 net426 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_96_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1320 total_design.core.regFile.register\[28\]\[23\] vssd1 vssd1 vccd1 vccd1 net2636
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout854_A _01947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10498__A0 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1331 total_design.core.regFile.register\[6\]\[31\] vssd1 vssd1 vccd1 vccd1 net2647
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08848_ _01746_ net537 vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__nand2_1
XANTENNA__10004__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1342 total_design.core.regFile.register\[4\]\[13\] vssd1 vssd1 vccd1 vccd1 net2658
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1353 total_design.core.regFile.register\[3\]\[10\] vssd1 vssd1 vccd1 vccd1 net2669
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1364 total_design.core.regFile.register\[15\]\[21\] vssd1 vssd1 vccd1 vccd1 net2680
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07902__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1375 total_design.core.regFile.register\[7\]\[15\] vssd1 vssd1 vccd1 vccd1 net2691
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1386 total_design.core.regFile.register\[7\]\[10\] vssd1 vssd1 vccd1 vccd1 net2702
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout642_X net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1397 total_design.core.regFile.register\[22\]\[12\] vssd1 vssd1 vccd1 vccd1 net2713
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08779_ _02718_ total_design.core.data_mem.data_cpu_i\[12\] vssd1 vssd1 vccd1 vccd1
+ _04034_ sky130_fd_sc_hd__and2b_1
XFILLER_0_68_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10810_ net518 _05049_ _05064_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_0_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11790_ net1787 net954 _05699_ _01793_ vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07115__B1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11998__B1 _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10741_ total_design.core.regFile.register\[0\]\[16\] net356 vssd1 vssd1 vccd1 vccd1
+ _01015_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout907_X net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13460_ clknet_leaf_143_clk _00927_ net1175 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10672_ net231 net1963 net361 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12411_ _01666_ _01667_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_11_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13391_ clknet_leaf_147_clk _00858_ net1152 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10674__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_20_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12342_ _01595_ _01598_ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__or2_1
XANTENNA__06453__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12273_ total_design.core.math.pc_val\[14\] total_design.core.program_count.imm_val_reg\[14\]
+ _06109_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06641__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14012_ clknet_leaf_98_clk _01192_ net1244 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11224_ _05362_ _05378_ _05482_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_31_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06929__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08394__A2 _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09591__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ _05405_ _05409_ _05413_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10262__X _05004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10106_ net209 net1932 net403 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__mux2_1
XANTENNA__12478__A1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13511__RESET_B net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11086_ _05327_ _05341_ _05344_ _05337_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_65_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_87_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08146__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10037_ net213 net2777 net410 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07354__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11988_ net531 _05842_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__nor2_4
XANTENNA__07106__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08303__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13727_ clknet_leaf_114_clk total_design.core.data_mem.stored_write_data\[2\] net1207
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[2\] sky130_fd_sc_hd__dfrtp_1
X_10939_ _05150_ _05168_ _05175_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_173_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13658_ clknet_leaf_55_clk total_design.core.data_mem.data_write_adr_i\[30\] net1114
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08843__A total_design.core.ctrl.instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12609_ clknet_leaf_122_clk _00076_ net1165 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10584__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13589_ clknet_leaf_34_clk total_design.core.data_mem.data_bus_i\[25\] net1066 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[25\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_11_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06632__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09820_ net283 net2329 net434 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__mux2_1
Xfanout407 net408 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_8
Xfanout418 net421 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_6
Xfanout429 _04977_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_129_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07593__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09751_ net268 net2391 net442 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__mux2_1
X_06963_ total_design.core.regFile.register\[29\]\[8\] net657 _02508_ _02512_ _02513_
+ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_78_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_33_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08702_ _00022_ _00021_ _00038_ _00037_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__or4_1
XANTENNA__08137__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09682_ net904 _04907_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__or2_1
X_06894_ _02448_ vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[7\] sky130_fd_sc_hd__inv_2
XANTENNA__07345__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ total_design.lcd_display.cnt_500hz\[11\] total_design.lcd_display.cnt_500hz\[10\]
+ total_design.lcd_display.cnt_500hz\[13\] total_design.lcd_display.cnt_500hz\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__or4_1
XANTENNA__08737__B _02845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08564_ total_design.data_in_BUS\[19\] net341 net718 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[19\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__06538__A _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07515_ net552 total_design.core.data_mem.data_cpu_i\[18\] total_design.core.ctrl.imm_32\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08495_ net933 total_design.keypad0.key_out\[10\] _03846_ vssd1 vssd1 vccd1 vccd1
+ _03847_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout435_A _04973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_138_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07446_ total_design.core.regFile.register\[1\]\[17\] net827 net790 total_design.core.regFile.register\[24\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__a22o_1
XANTENNA__06856__C1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10494__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout602_A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07377_ total_design.core.regFile.register\[22\]\[16\] net675 net626 total_design.core.regFile.register\[14\]\[16\]
+ _02903_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__a221o_1
XANTENNA__06871__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06544__Y _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07369__A total_design.core.ctrl.instruction\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09116_ _04126_ _04365_ net326 vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__mux2_1
X_06328_ net997 net1266 _01905_ _01906_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06623__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09047_ net466 _04169_ _04298_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__o21a_1
X_06259_ total_design.core.data_adr_o\[27\] _01837_ net962 vssd1 vssd1 vccd1 vccd1
+ _01838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold450 total_design.lcd_display.row_2\[119\] vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold461 total_design.lcd_display.row_2\[53\] vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout971_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap180 _05316_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_1
Xhold472 total_design.lcd_display.row_1\[24\] vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_147_Left_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09573__A1 total_design.core.data_cpu_o\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11619__A _05478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold483 total_design.core.mem_ctrl.state\[2\] vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 net101 vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07584__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout930 _01807_ vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_4
Xfanout941 _03675_ vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06212__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09949_ net163 net2291 net423 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__mux2_1
Xfanout952 _01914_ vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__buf_2
Xfanout963 _01770_ vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_69_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout857_X net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08128__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout974 net975 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__clkbuf_2
Xfanout985 total_design.core.disable_pc vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_4
Xfanout996 total_design.core.program_count.ALU_out_reg vssd1 vssd1 vccd1 vccd1 net996
+ sky130_fd_sc_hd__clkbuf_2
X_12960_ clknet_leaf_2_clk _00427_ net1011 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 net122 vssd1 vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07336__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11911_ _03982_ _05774_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__nor2_1
Xhold1161 total_design.data_in_BUS\[24\] vssd1 vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 total_design.core.regFile.register\[23\]\[18\] vssd1 vssd1 vccd1 vccd1 net2488
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10669__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12891_ clknet_leaf_144_clk _00358_ net1174 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1183 total_design.core.regFile.register\[11\]\[6\] vssd1 vssd1 vccd1 vccd1 net2499
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 total_design.core.regFile.register\[8\]\[19\] vssd1 vssd1 vccd1 vccd1 net2510
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14199__RESET_B net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11842_ _01724_ total_design.lcd_display.currentState\[1\] total_design.lcd_display.currentState\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_156_Left_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08366__C _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14561_ net1281 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
X_11773_ net1720 net955 net301 _01789_ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08934__Y _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13512_ clknet_leaf_172_clk _00979_ net1056 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10724_ total_design.core.instr_fetch net507 vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__or2_4
XFILLER_0_32_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14492_ clknet_leaf_27_clk _01559_ net1074 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_71_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13443_ clknet_leaf_16_clk _00910_ net1024 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11801__B net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10655_ net169 net2297 net476 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__mux2_1
XANTENNA__06862__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12185__A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11520__C _05479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13374_ clknet_leaf_175_clk _00841_ net1053 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload17 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__bufinv_16
Xclkload28 clknet_leaf_181_clk vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__bufinv_16
X_10586_ net181 net2204 net371 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload39 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__clkinv_4
X_12325_ net990 _04737_ net894 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12148__B1 _05971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_165_Left_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12256_ total_design.core.math.pc_val\[12\] total_design.core.program_count.imm_val_reg\[12\]
+ _06094_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11207_ _05450_ _05455_ _05465_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_121_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07726__B _03234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09564__B2 _04443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12187_ total_design.core.math.pc_val\[5\] total_design.core.program_count.imm_val_reg\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__or2_1
XANTENNA__11371__A1 total_design.core.data_bus_o\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11138_ _05382_ _05383_ _05396_ _05386_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__o31a_1
XANTENNA__11108__D1 _05028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08119__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ net351 _05281_ _05285_ _05290_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__nand4_1
Xclkbuf_leaf_0_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10579__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5__f_clk_X clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07300_ total_design.core.regFile.register\[5\]\[14\] net809 net764 total_design.core.regFile.register\[6\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__a22o_1
XANTENNA__06508__D net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08280_ net1357 net557 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[30\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07231_ total_design.core.regFile.register\[31\]\[13\] net601 _02752_ _02766_ vssd1
+ vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__a211o_1
XANTENNA__06853__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09388__B net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07162_ total_design.core.regFile.register\[19\]\[12\] net641 net568 total_design.core.regFile.register\[12\]\[12\]
+ _02700_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07093_ _02634_ _02636_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__nand2_2
XANTENNA__06605__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout204 _04760_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_2
Xfanout215 _04681_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_2
Xfanout226 net227 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__dlymetal6s2s_1
X_09803_ net198 net2834 net439 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__mux2_1
Xfanout237 net239 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_1
XANTENNA__07030__A2 _01994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07995_ total_design.core.regFile.register\[29\]\[28\] net656 net574 total_design.core.regFile.register\[24\]\[28\]
+ _03491_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__a221o_1
Xfanout259 net260 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout385_A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _04956_ _04321_ net329 _04877_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__o2bb2a_1
X_06946_ total_design.core.regFile.register\[18\]\[8\] net610 net603 total_design.core.regFile.register\[31\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09665_ _03459_ _03461_ _04872_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10489__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06877_ total_design.core.regFile.register\[13\]\[6\] net788 net778 total_design.core.regFile.register\[22\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout552_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13804__D total_design.core.data_mem.data_cpu_i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08616_ total_design.keypad0.next_rows\[1\] total_design.keypad0.next_rows\[3\] total_design.keypad0.next_rows\[2\]
+ vssd1 vssd1 vccd1 vccd1 total_design.keypad0.next_rows\[0\] sky130_fd_sc_hd__nand3_1
XFILLER_0_96_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09596_ _04807_ _04823_ _03373_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__o21a_1
X_08547_ net717 _03895_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[11\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout817_A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12090__A2 _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ _03827_ _03829_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07429_ total_design.core.regFile.register\[26\]\[17\] net644 net573 total_design.core.regFile.register\[24\]\[17\]
+ _02951_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__a221o_1
XFILLER_0_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06844__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout605_X net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10440_ net239 net2809 net382 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08949__D_N total_design.core.ctrl.instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10371_ net249 net2040 net487 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__mux2_1
X_12110_ total_design.lcd_display.row_1\[69\] _05804_ _05829_ total_design.lcd_display.row_1\[109\]
+ _05966_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__a221o_1
X_13090_ clknet_leaf_129_clk _00557_ net1193 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_148_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12041_ total_design.lcd_display.row_2\[90\] _05837_ _05845_ total_design.lcd_display.row_2\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__a22o_1
Xhold280 total_design.lcd_display.row_2\[7\] vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 total_design.lcd_display.row_1\[76\] vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07557__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07021__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout760 net762 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__clkbuf_8
Xfanout771 net772 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__buf_4
Xfanout782 _01988_ vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__buf_4
X_13992_ clknet_leaf_73_clk _01172_ net1221 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_184_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout793 _01982_ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__buf_4
XFILLER_0_172_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_161_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ clknet_leaf_160_clk _00410_ net1150 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10399__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12874_ clknet_leaf_22_clk _00341_ net1049 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11825_ total_design.lcd_display.cnt_20ms\[13\] _05713_ net1879 vssd1 vssd1 vccd1
+ vccd1 _05716_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_199_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11371__X _05630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14544_ net1316 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XFILLER_0_134_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11756_ net1743 net959 net292 total_design.core.data_bus_o\[28\] vssd1 vssd1 vccd1
+ vccd1 _01384_ sky130_fd_sc_hd__a22o_1
XANTENNA__12081__A2 _05834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08393__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ net224 net1976 net360 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__mux2_1
X_14475_ clknet_leaf_39_clk _01542_ net1091 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_11687_ total_design.bus_full wishbone.prev_BUSY_O net935 vssd1 vssd1 vccd1 vccd1
+ _05690_ sky130_fd_sc_hd__and3b_1
XFILLER_0_126_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_122_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13426_ clknet_leaf_145_clk _00893_ net1177 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10638_ net237 net2405 net479 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__mux2_1
XANTENNA__09001__B _03112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload106 clknet_leaf_160_clk vssd1 vssd1 vccd1 vccd1 clkload106/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload117 clknet_leaf_167_clk vssd1 vssd1 vccd1 vccd1 clkload117/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload128 clknet_leaf_143_clk vssd1 vssd1 vccd1 vccd1 clkload128/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__06344__C total_design.core.ctrl.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_141_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload139 clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 clkload139/Y sky130_fd_sc_hd__clkinv_4
X_13357_ clknet_leaf_3_clk _00824_ net1013 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10569_ net249 net2403 net372 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12308_ _01573_ _01575_ _01576_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13288_ clknet_leaf_117_clk _00755_ net1162 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_137_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12239_ total_design.core.math.pc_val\[11\] total_design.core.program_count.imm_val_reg\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__nand2_1
XANTENNA__07548__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07012__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06800_ total_design.core.regFile.register\[25\]\[5\] net649 net629 total_design.core.regFile.register\[5\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__a22o_1
X_07780_ total_design.core.regFile.register\[29\]\[24\] net799 net777 total_design.core.regFile.register\[22\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07472__A total_design.core.ctrl.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_06731_ total_design.core.regFile.register\[15\]\[4\] net846 net823 total_design.core.regFile.register\[19\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09450_ _04191_ _04303_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06662_ total_design.core.regFile.register\[13\]\[2\] net667 net563 total_design.core.regFile.register\[3\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__a22o_1
XANTENNA__10102__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08401_ _03755_ _03756_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06519__C net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09381_ _02893_ net701 _04619_ net533 vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a211o_1
X_06593_ total_design.core.regFile.register\[20\]\[1\] net746 net739 net735 vssd1
+ vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__and4_1
XFILLER_0_15_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10607__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ net1454 net938 _03700_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[23\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09399__A _02868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07079__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06375__X _01951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08734__C _02492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08263_ net1416 net559 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[13\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__06826__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13710__Q total_design.core.data_cpu_o\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout133_A _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06535__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07214_ net550 _02749_ _02750_ vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[13\]
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_27_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08194_ _03647_ _03648_ _03649_ _03650_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07145_ net300 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[11\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_30_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1042_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07787__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07076_ total_design.core.regFile.register\[27\]\[10\] net779 _02620_ vssd1 vssd1
+ vccd1 vccd1 _02621_ sky130_fd_sc_hd__a21o_1
XANTENNA__07251__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07539__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12532__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07003__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout767_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10801__A total_design.core.data_bus_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ total_design.core.regFile.register\[31\]\[28\] net833 net803 total_design.core.regFile.register\[8\]\[28\]
+ _03475_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09717_ net315 _04193_ _04770_ _04940_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__a31o_1
X_06929_ total_design.core.regFile.register\[5\]\[7\] net809 net779 total_design.core.regFile.register\[27\]\[7\]
+ _02470_ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout934_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10012__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ _04269_ _04271_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__nor2_1
XFILLER_0_167_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07711__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09801__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09579_ _03329_ net705 _04806_ _04808_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__a22o_1
X_11610_ _05628_ net1762 net140 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12063__A2 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12590_ clknet_leaf_188_clk _00057_ net1028 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11541_ net1511 _05636_ net146 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06817__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14260_ clknet_leaf_102_clk _01439_ net1239 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.currentState\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_11472_ net1522 _05657_ net153 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__mux2_1
XANTENNA__07490__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire457 _03131_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_4
X_13211_ clknet_leaf_150_clk _00678_ net1147 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10423_ net174 net2055 net386 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__mux2_1
X_14191_ clknet_leaf_80_clk _01371_ net1221 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10682__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07778__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13142_ clknet_leaf_152_clk _00609_ net1138 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10354_ net187 net2617 net489 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__mux2_1
XANTENNA__07242__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06450__B1 _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ clknet_leaf_150_clk _00540_ net1145 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10285_ net200 net2801 net498 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_163_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12024_ total_design.lcd_display.row_1\[97\] _05810_ _05821_ total_design.lcd_display.row_1\[41\]
+ _05884_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_163_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_168_Right_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06202__A0 total_design.core.instr_mem.instruction_adr_i\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08742__A2 _03602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07950__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 net592 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__buf_4
XFILLER_0_73_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13975_ clknet_leaf_84_clk _01155_ net1243 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_12926_ clknet_leaf_181_clk _00393_ net1140 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07702__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12857_ clknet_leaf_195_clk _00324_ net1012 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11808_ _05705_ _05706_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__and2b_1
XANTENNA__12054__A2 _05832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12788_ clknet_leaf_142_clk _00255_ net1175 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06636__A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11739_ net1744 net958 net290 total_design.core.data_bus_o\[11\] vssd1 vssd1 vccd1
+ vccd1 _01367_ sky130_fd_sc_hd__a22o_1
X_14527_ net1299 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XANTENNA__06808__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09207__B1 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14458_ clknet_leaf_53_clk net1499 net1095 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07481__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ clknet_leaf_123_clk _00876_ net1188 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14389_ clknet_leaf_136_clk _01530_ net1180 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06642__Y total_design.core.data_mem.data_cpu_i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07233__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08950_ _01922_ _02445_ _04202_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__nor3_1
XANTENNA__12514__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09682__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07901_ total_design.core.regFile.register\[23\]\[26\] net679 net646 total_design.core.regFile.register\[26\]\[26\]
+ _03401_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__a221o_1
XANTENNA__06521__D net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08881_ _04131_ _04134_ net459 vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_102_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07832_ total_design.core.regFile.register\[17\]\[25\] net820 _03333_ _03335_ vssd1
+ vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__a211o_1
X_07763_ total_design.core.regFile.register\[21\]\[23\] net597 net566 total_design.core.regFile.register\[12\]\[23\]
+ _03256_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__a221o_1
X_09502_ total_design.core.math.pc_val\[20\] _04715_ vssd1 vssd1 vccd1 vccd1 _04736_
+ sky130_fd_sc_hd__nor2_1
X_06714_ total_design.core.regFile.register\[30\]\[3\] net659 net632 total_design.core.regFile.register\[16\]\[3\]
+ _02278_ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07694_ _03197_ _03199_ _03201_ _03203_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__or4_1
XFILLER_0_116_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ _04573_ _04669_ net328 vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__mux2_1
XANTENNA__11723__Y _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06645_ _02116_ _02187_ _02185_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09364_ net314 _04408_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__or2_2
XFILLER_0_136_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12045__A2 _05819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06576_ _02142_ _02144_ _02148_ net874 total_design.core.regFile.register\[0\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[1\] sky130_fd_sc_hd__o32a_4
XPHY_EDGE_ROW_111_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08315_ total_design.core.data_mem.data_write_adr_reg\[15\] net548 net540 total_design.core.data_mem.data_read_adr_reg\[15\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_23_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09295_ _04525_ _04537_ _04124_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_43_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout515_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1257_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08246_ net1395 net543 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[29\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_16_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11598__S net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08177_ net890 _03138_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[20\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1045_X net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07128_ total_design.core.regFile.register\[10\]\[11\] net837 _02668_ _02669_ vssd1
+ vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_132_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07224__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07059_ total_design.core.regFile.register\[7\]\[10\] net651 net632 total_design.core.regFile.register\[16\]\[10\]
+ _02603_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a221o_1
XANTENNA__10007__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1212_X net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10070_ net220 net2347 net407 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07932__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06220__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13760_ clknet_leaf_61_clk total_design.core.data_mem.stored_data_adr\[3\] net1216
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[3\] sky130_fd_sc_hd__dfrtp_1
X_10972_ _05217_ _05225_ _05227_ _05229_ _05230_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_67_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12711_ clknet_leaf_19_clk _00178_ net1049 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13691_ clknet_leaf_55_clk total_design.core.data_mem.data_read_adr_i\[31\] net1113
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[31\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10677__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07160__A1 total_design.core.ctrl.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06727__Y _02292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12642_ clknet_leaf_129_clk _00109_ net1193 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12036__A2 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12573_ clknet_leaf_9_clk _00040_ net1020 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07999__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14312_ clknet_leaf_63_clk _01473_ net1124 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_11524_ net1591 _05635_ net147 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__mux2_1
X_14243_ clknet_leaf_109_clk _01423_ net1228 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11455_ net1569 _05477_ net155 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__mux2_1
XANTENNA__09486__B _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11547__A1 _05645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ net242 net2385 net385 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__mux2_1
X_14174_ clknet_leaf_60_clk _01354_ net1132 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06191__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11386_ _05584_ _05642_ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__o21a_2
XFILLER_0_22_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13125_ clknet_leaf_117_clk _00592_ net1212 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10337_ net263 net2827 net490 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13056_ clknet_leaf_3_clk _00523_ net1013 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10268_ net259 net2174 net499 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__mux2_1
X_12007_ total_design.lcd_display.row_1\[64\] _05804_ _05810_ total_design.lcd_display.row_1\[96\]
+ _05828_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10199_ _04474_ net392 _04996_ vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07923__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09007__A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13958_ clknet_leaf_101_clk _01138_ net1237 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08846__A total_design.core.ctrl.instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_159_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12909_ clknet_leaf_6_clk _00376_ net1016 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10587__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13889_ clknet_leaf_96_clk _01069_ net1254 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06430_ _02001_ _02002_ _02003_ _02005_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__or4_1
XFILLER_0_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12027__A2 _05838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06366__A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09428__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06361_ net951 net950 _01738_ net965 net952 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08100__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11786__A1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08100_ total_design.core.regFile.register\[10\]\[30\] net618 net610 total_design.core.regFile.register\[18\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09080_ _04213_ _04330_ net461 vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__mux2_1
X_06292_ _01859_ _01861_ _01866_ _01868_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__and4_1
XANTENNA__07454__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08031_ total_design.core.regFile.register\[5\]\[29\] net806 _01992_ total_design.core.regFile.register\[20\]\[29\]
+ _03514_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06662__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold802 total_design.core.regFile.register\[27\]\[23\] vssd1 vssd1 vccd1 vccd1 net2118
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold813 total_design.core.regFile.register\[10\]\[18\] vssd1 vssd1 vccd1 vccd1 net2129
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 total_design.core.regFile.register\[6\]\[20\] vssd1 vssd1 vccd1 vccd1 net2140
+ sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap532 _05001_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_4
XFILLER_0_101_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold835 total_design.core.regFile.register\[29\]\[14\] vssd1 vssd1 vccd1 vccd1 net2151
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 total_design.core.regFile.register\[22\]\[17\] vssd1 vssd1 vccd1 vccd1 net2162
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold857 total_design.core.regFile.register\[20\]\[19\] vssd1 vssd1 vccd1 vccd1 net2173
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09683__Y _04909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09982_ net165 net2847 net420 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__mux2_1
Xhold868 total_design.data_in_BUS\[25\] vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 total_design.core.regFile.register\[16\]\[20\] vssd1 vssd1 vccd1 vccd1 net2195
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08933_ net969 net537 vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1502 total_design.core.regFile.register\[20\]\[10\] vssd1 vssd1 vccd1 vccd1 net2818
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08864_ total_design.core.ctrl.instruction\[7\] total_design.core.ctrl.instruction\[8\]
+ net556 vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__o21a_1
Xhold1513 total_design.core.regFile.register\[17\]\[4\] vssd1 vssd1 vccd1 vccd1 net2829
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1005_A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1524 total_design.core.regFile.register\[23\]\[0\] vssd1 vssd1 vccd1 vccd1 net2840
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07914__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1535 total_design.core.regFile.register\[18\]\[7\] vssd1 vssd1 vccd1 vccd1 net2851
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07815_ total_design.core.regFile.register\[4\]\[24\] net621 net583 total_design.core.regFile.register\[6\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__a22o_1
XANTENNA__11166__B _05184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1546 total_design.core.regFile.register\[6\]\[19\] vssd1 vssd1 vccd1 vccd1 net2862
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08795_ _04045_ _04046_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__nand2b_1
Xhold1557 total_design.core.regFile.register\[16\]\[8\] vssd1 vssd1 vccd1 vccd1 net2873
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1568 total_design.data_in_BUS\[25\] vssd1 vssd1 vccd1 vccd1 net2884 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_88_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07746_ _03253_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[23\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__08756__A _03253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09204__X _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ net749 _03187_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[21\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10497__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout632_A _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ net904 _04653_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06628_ total_design.core.regFile.register\[16\]\[2\] net854 net775 total_design.core.regFile.register\[22\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__a22o_1
XANTENNA__12018__A2 _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07693__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06350__C1 _01915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14266__Q total_design.core.math.pc_val\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09347_ _04587_ _04586_ _04582_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__or3b_2
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06559_ total_design.core.regFile.register\[14\]\[1\] net920 net916 net946 vssd1
+ vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09278_ _02613_ _02633_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08229_ net1461 net544 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[12\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__06653__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07819__B _03322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11529__A1 _05663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11240_ _05490_ _05493_ _05496_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__a21oi_2
XANTENNA__06215__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10201__A1 _04495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ _05425_ _05429_ _05422_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__o21ai_1
X_10122_ net244 net2686 net398 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__mux2_1
XANTENNA__09355__C1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ _04115_ _04986_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__nand2_1
XANTENNA__07905__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ clknet_leaf_113_clk total_design.core.data_mem.data_cpu_i\[21\] net1203 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[21\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09658__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10955_ _05197_ _05203_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__and2b_1
X_13743_ clknet_leaf_72_clk total_design.core.data_mem.stored_write_data\[18\] net1205
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[18\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_27_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13674_ clknet_leaf_55_clk total_design.core.data_mem.data_read_adr_i\[14\] net1120
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[14\] sky130_fd_sc_hd__dfrtp_1
X_10886_ _05143_ _05144_ _05127_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__a21oi_4
XANTENNA__07684__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14176__Q net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12625_ clknet_leaf_151_clk _00092_ net1145 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12556_ net1414 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07436__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09830__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11507_ net1576 _05652_ net151 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12487_ net979 total_design.core.instr_mem.instruction_i\[7\] vssd1 vssd1 vccd1 vccd1
+ _01698_ sky130_fd_sc_hd__and2b_1
Xhold109 total_design.core.instr_mem.instruction_adr_stored\[27\] vssd1 vssd1 vccd1
+ vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
X_14226_ clknet_leaf_57_clk _01406_ net1118 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dfrtp_1
X_11438_ net1803 _05671_ net157 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__mux2_1
XANTENNA_output94_A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14157_ clknet_leaf_31_clk _01337_ net1060 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08936__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11369_ total_design.core.data_bus_o\[23\] net699 net511 vssd1 vssd1 vccd1 vccd1
+ _05628_ sky130_fd_sc_hd__a21o_2
XFILLER_0_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13108_ clknet_leaf_141_clk _00575_ net1182 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14088_ clknet_leaf_110_clk _01268_ net1227 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08149__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13039_ clknet_leaf_161_clk _00506_ net1151 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12496__A2 total_design.core.ctrl.instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_119_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1160 net1162 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__clkbuf_4
Xfanout1171 net1172 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__clkbuf_4
Xfanout1182 net1201 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11417__D _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1193 net1194 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__clkbuf_4
X_07600_ total_design.core.regFile.register\[15\]\[20\] net846 net827 total_design.core.regFile.register\[1\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__a22o_1
XANTENNA__08847__Y _04102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08580_ _03723_ net880 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[1\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07531_ total_design.core.regFile.register\[21\]\[19\] net598 net590 total_design.core.regFile.register\[1\]\[19\]
+ _03047_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10110__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07462_ total_design.core.regFile.register\[2\]\[17\] net783 _01992_ total_design.core.regFile.register\[20\]\[17\]
+ _02985_ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_83_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08863__X _04117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09201_ total_design.core.math.pc_val\[5\] total_design.core.math.pc_val\[6\] total_design.core.math.pc_val\[7\]
+ _04371_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__and4_1
XFILLER_0_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06413_ total_design.core.regFile.register\[27\]\[0\] net928 net915 net912 vssd1
+ vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__and4_1
XFILLER_0_91_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07393_ total_design.core.regFile.register\[12\]\[16\] _01994_ _01995_ total_design.core.regFile.register\[28\]\[16\]
+ _02919_ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__a221o_1
XFILLER_0_162_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11759__A1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09132_ net323 _04230_ net314 vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__a21o_1
XANTENNA__11759__B2 total_design.core.data_bus_o\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06344_ net971 net973 total_design.core.ctrl.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ _01920_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_174_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07427__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06383__X _01959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09063_ _04313_ _04314_ net452 vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_5_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06635__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06275_ total_design.core.data_adr_o\[2\] _01853_ net963 vssd1 vssd1 vccd1 vccd1
+ _01854_ sky130_fd_sc_hd__mux2_2
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08014_ _03464_ _03466_ _03509_ _03463_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_142_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold610 total_design.core.regFile.register\[14\]\[23\] vssd1 vssd1 vccd1 vccd1 net1926
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 total_design.core.regFile.register\[8\]\[2\] vssd1 vssd1 vccd1 vccd1 net1937
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold632 total_design.core.regFile.register\[2\]\[7\] vssd1 vssd1 vccd1 vccd1 net1948
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 total_design.core.regFile.register\[2\]\[26\] vssd1 vssd1 vccd1 vccd1 net1959
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 total_design.core.regFile.register\[24\]\[25\] vssd1 vssd1 vccd1 vccd1 net1970
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 total_design.core.regFile.register\[3\]\[13\] vssd1 vssd1 vccd1 vccd1 net1981
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 total_design.core.regFile.register\[14\]\[26\] vssd1 vssd1 vccd1 vccd1 net1992
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold687 total_design.core.regFile.register\[22\]\[20\] vssd1 vssd1 vccd1 vccd1 net2003
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07060__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold698 total_design.core.regFile.register\[0\]\[21\] vssd1 vssd1 vccd1 vccd1 net2014
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ net230 net2190 net421 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout582_A _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13807__D total_design.core.data_mem.data_cpu_i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08916_ _04167_ _04169_ net465 vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__mux2_1
XANTENNA__09888__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09896_ net238 net2823 net427 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__mux2_1
Xhold1310 total_design.core.regFile.register\[19\]\[18\] vssd1 vssd1 vccd1 vccd1 net2626
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1321 total_design.core.regFile.register\[4\]\[9\] vssd1 vssd1 vccd1 vccd1 net2637
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11695__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1332 total_design.core.regFile.register\[18\]\[10\] vssd1 vssd1 vccd1 vccd1 net2648
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1343 total_design.core.regFile.register\[22\]\[25\] vssd1 vssd1 vccd1 vccd1 net2659
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ net968 _04101_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__nor2_2
Xhold1354 total_design.core.regFile.register\[13\]\[26\] vssd1 vssd1 vccd1 vccd1 net2670
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout847_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1365 total_design.core.regFile.register\[5\]\[17\] vssd1 vssd1 vccd1 vccd1 net2681
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1376 total_design.core.regFile.register\[18\]\[22\] vssd1 vssd1 vccd1 vccd1 net2692
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1387 total_design.core.regFile.register\[26\]\[21\] vssd1 vssd1 vccd1 vccd1 net2703
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08778_ _04005_ _04015_ _04032_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__or3_1
Xhold1398 total_design.core.regFile.register\[12\]\[13\] vssd1 vssd1 vccd1 vccd1 net2714
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07729_ total_design.core.regFile.register\[14\]\[23\] net861 net767 total_design.core.regFile.register\[7\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10020__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10740_ total_design.core.regFile.register\[0\]\[15\] net356 vssd1 vssd1 vccd1 vccd1
+ _01014_ sky130_fd_sc_hd__and2_1
XANTENNA__07666__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06874__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10671_ net236 net2004 net363 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12410_ total_design.core.math.pc_val\[29\] net989 _01666_ vssd1 vssd1 vccd1 vccd1
+ _01668_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08933__B net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13390_ clknet_leaf_189_clk _00857_ net1029 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12341_ _01604_ _01605_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08091__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06453__B _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12272_ total_design.core.math.pc_val\[14\] net527 _06106_ _06112_ vssd1 vssd1 vccd1
+ vccd1 _01484_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14011_ clknet_leaf_94_clk _01191_ net1257 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11223_ _05372_ _05378_ _05362_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__and3b_1
XANTENNA__10690__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09040__A1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07051__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ _05399_ _05406_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_105_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10105_ net218 net2626 net402 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__mux2_1
X_11085_ _05342_ _05343_ net351 _05272_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__o2bb2a_1
X_10036_ net220 net2343 net412 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__mux2_1
XANTENNA__11374__X _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08303__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11987_ net531 _05800_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__nor2_4
XANTENNA__09004__B net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13726_ clknet_leaf_112_clk total_design.core.data_mem.stored_write_data\[1\] net1207
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[1\] sky130_fd_sc_hd__dfrtp_1
X_10938_ _05195_ _05196_ _05180_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07657__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13657_ clknet_leaf_54_clk total_design.core.data_mem.data_write_adr_i\[29\] net1113
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[29\] sky130_fd_sc_hd__dfrtp_1
X_10869_ _05113_ _05117_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__nor2_1
XANTENNA__08843__B _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12608_ clknet_leaf_2_clk _00075_ net1011 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13588_ clknet_leaf_33_clk total_design.core.data_mem.data_bus_i\[24\] net1070 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11610__A0 _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08562__C net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12539_ total_design.core.ctrl.instruction\[31\] net885 _02149_ _03091_ net550 vssd1
+ vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[23\] sky130_fd_sc_hd__a221o_1
XANTENNA__08082__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07290__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12166__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14209_ clknet_leaf_60_clk _01389_ net1131 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout408 net409 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_8
Xfanout419 net421 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_6
XANTENNA__10105__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ net279 total_design.core.regFile.register\[29\]\[2\] net442 vssd1 vssd1 vccd1
+ vccd1 _00073_ sky130_fd_sc_hd__mux2_1
X_06962_ total_design.core.regFile.register\[7\]\[8\] net654 net591 total_design.core.regFile.register\[1\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a22o_1
X_08701_ net1783 _03953_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__xor2_1
XANTENNA__11677__A0 _05648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09681_ _04905_ _04906_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_33_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06893_ net721 _02446_ _02447_ _02444_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__o211a_2
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08632_ _03921_ net711 _03920_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_85_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07896__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08737__C _02893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08563_ net1946 net339 net718 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[18\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_81_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07514_ total_design.core.regFile.register\[0\]\[18\] net873 _03028_ _03034_ vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[18\] sky130_fd_sc_hd__o22a_4
XFILLER_0_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08494_ net933 total_design.keypad0.key_out\[10\] _03810_ vssd1 vssd1 vccd1 vccd1
+ _03846_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07648__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07445_ _02968_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1072_A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07376_ total_design.core.regFile.register\[5\]\[16\] net629 net586 total_design.core.regFile.register\[28\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11601__A0 _05655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09115_ net460 _04364_ _04363_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__a21oi_1
X_06327_ _01766_ _01768_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06608__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08073__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07281__B1 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09046_ net465 _04175_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__nand2_1
X_06258_ total_design.core.instr_mem.instruction_adr_i\[27\] total_design.core.instr_mem.instruction_adr_stored\[27\]
+ net981 vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06841__X total_design.core.ctrl.imm_32\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09558__C1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold440 total_design.lcd_display.row_1\[98\] vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06189_ _01767_ _01768_ _01769_ _01761_ vssd1 vssd1 vccd1 vccd1 total_design.core.mem_ctrl.next_state\[0\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10804__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold451 net60 vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold462 net48 vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 total_design.lcd_display.row_2\[30\] vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07033__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09573__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold484 total_design.lcd_display.row_2\[26\] vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 _01362_ vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout964_A _01770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout585_X net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout920 net924 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_2
Xfanout931 total_design.keypad0.key_out\[14\] vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_2
Xfanout942 _03674_ vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__buf_2
XANTENNA__10015__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ net165 total_design.core.regFile.register\[24\]\[30\] net424 vssd1 vssd1
+ vccd1 vccd1 _00261_ sky130_fd_sc_hd__mux2_1
Xfanout953 _01911_ vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__buf_2
Xfanout964 _01770_ vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11668__A0 _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout975 net978 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__buf_2
XANTENNA__09804__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout986 total_design.keypad0.key_clk vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout997 total_design.core.data_mem.data_write vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ net169 net2280 net430 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 total_design.core.regFile.register\[1\]\[11\] vssd1 vssd1 vccd1 vccd1 net2456
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 total_design.core.regFile.register\[14\]\[13\] vssd1 vssd1 vccd1 vccd1 net2467
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ net999 _05778_ _05786_ _03907_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__o22a_1
Xhold1162 total_design.core.regFile.register\[19\]\[5\] vssd1 vssd1 vccd1 vccd1 net2478
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07391__Y _02918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1173 total_design.core.regFile.register\[30\]\[29\] vssd1 vssd1 vccd1 vccd1 net2489
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07887__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12890_ clknet_leaf_133_clk _00357_ net1196 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 total_design.core.regFile.register\[10\]\[3\] vssd1 vssd1 vccd1 vccd1 net2500
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1195 total_design.core.regFile.register\[21\]\[2\] vssd1 vssd1 vccd1 vccd1 net2511
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11841_ total_design.lcd_display.currentState\[4\] total_design.lcd_display.currentState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_16_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14560_ net1280 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
X_11772_ net1798 net955 net301 _01800_ vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07639__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10723_ net162 net2359 net360 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__mux2_1
X_13511_ clknet_leaf_174_clk _00978_ net1058 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06847__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10685__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14491_ clknet_leaf_37_clk _01558_ net1076 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10654_ net172 net2187 net478 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__mux2_1
X_13442_ clknet_leaf_126_clk _00909_ net1193 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12185__B _02395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14454__Q total_design.core.instr_mem.instruction_adr_i\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13373_ clknet_leaf_14_clk _00840_ net1026 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10585_ net185 net2160 net371 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__mux2_1
XANTENNA__11520__D _05675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload18 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload18/X sky130_fd_sc_hd__clkbuf_8
Xclkload29 clknet_leaf_183_clk vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__clkinvlp_4
X_12324_ _01588_ _01589_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_118_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07272__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07811__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11369__X _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12255_ total_design.core.math.pc_val\[12\] net527 _06090_ _06097_ vssd1 vssd1 vccd1
+ vccd1 _01482_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11206_ _05445_ _05464_ _05447_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07024__B1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12186_ total_design.core.math.pc_val\[4\] total_design.core.program_count.imm_val_reg\[4\]
+ _06030_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11371__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ _05384_ _05388_ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__nor2_1
XANTENNA__11659__A0 _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09316__A2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ _05286_ _05290_ _05326_ _05184_ _05045_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__a32o_1
X_10019_ _04115_ _04984_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__nand2_1
XANTENNA__10331__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07878__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12084__B1 _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13709_ clknet_leaf_27_clk total_design.core.data_mem.stored_read_data\[16\] net1073
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[16\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10595__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06645__Y _02213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07230_ total_design.core.regFile.register\[22\]\[13\] net674 _02764_ _02765_ vssd1
+ vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__a211o_1
XFILLER_0_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07161_ total_design.core.regFile.register\[9\]\[12\] net665 net598 total_design.core.regFile.register\[21\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07092_ _02613_ _02633_ vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07802__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout205 _04740_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_2
Xfanout216 _04699_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_2
X_09802_ net202 net2871 net439 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__mux2_1
Xfanout227 _04636_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_2
Xfanout238 net239 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
X_07994_ total_design.core.regFile.register\[22\]\[28\] net675 net586 total_design.core.regFile.register\[28\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__a22o_1
Xfanout249 net252 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_52_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06945_ _02449_ _02490_ _02489_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__a21boi_2
X_09733_ net467 _04918_ _04955_ net330 vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout280_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07318__A1 total_design.core.ctrl.instruction\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout378_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10322__A0 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ net177 net2393 net455 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__mux2_1
X_06876_ total_design.core.regFile.register\[14\]\[6\] net863 _02432_ vssd1 vssd1
+ vccd1 vccd1 _02433_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08615_ _03908_ vssd1 vssd1 vccd1 vccd1 total_design.keypad0.next_rows\[2\] sky130_fd_sc_hd__inv_2
X_09595_ _03373_ _04807_ _04823_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__nor3_1
XFILLER_0_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12075__B1 _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08546_ net2880 net342 _03894_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06836__X _02395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08477_ _03827_ _03829_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout712_A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1075_X net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07428_ total_design.core.regFile.register\[19\]\[17\] net640 net620 total_design.core.regFile.register\[4\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07359_ _02871_ _02874_ _02888_ net876 total_design.core.regFile.register\[0\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[15\] sky130_fd_sc_hd__o32a_4
XFILLER_0_165_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08046__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10370_ net264 net2353 net487 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10805__Y _05064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09029_ net245 net1889 net454 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12040_ total_design.lcd_display.row_1\[50\] _05840_ _05850_ total_design.lcd_display.row_2\[2\]
+ _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__a221o_1
XANTENNA__07006__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold270 total_design.lcd_display.row_1\[45\] vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06223__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold281 total_design.lcd_display.row_2\[121\] vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 total_design.lcd_display.row_1\[74\] vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10561__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout750 net753 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_2
Xfanout761 net762 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_8
Xfanout772 _01995_ vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_6
X_13991_ clknet_leaf_82_clk _01171_ net1241 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout783 _01986_ vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__clkbuf_8
Xfanout794 net797 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ clknet_leaf_189_clk _00409_ net1029 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_161_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ clknet_leaf_178_clk _00340_ net1033 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06532__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12066__B1 _05848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11824_ total_design.lcd_display.cnt_20ms\[13\] total_design.lcd_display.cnt_20ms\[14\]
+ _05713_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14543_ net1315 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
X_11755_ net1587 net958 net291 total_design.core.data_bus_o\[27\] vssd1 vssd1 vccd1
+ vccd1 _01383_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10706_ net232 net2664 net358 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14474_ clknet_leaf_40_clk _01541_ net1092 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11686_ wishbone.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13425_ clknet_leaf_148_clk _00892_ net1149 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10637_ net240 net2622 net479 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__mux2_1
Xclkload107 clknet_leaf_161_clk vssd1 vssd1 vccd1 vccd1 clkload107/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload118 clknet_leaf_168_clk vssd1 vssd1 vccd1 vccd1 clkload118/Y sky130_fd_sc_hd__inv_8
Xclkload129 clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 clkload129/Y sky130_fd_sc_hd__inv_6
XANTENNA__07245__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13356_ clknet_leaf_165_clk _00823_ net1158 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10568_ net264 net2767 net371 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06599__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_168_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11099__X _05358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12307_ _01573_ _01575_ net990 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13287_ clknet_leaf_176_clk _00754_ net1052 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10499_ net258 net2431 net483 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_15_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12238_ total_design.core.math.pc_val\[10\] total_design.core.program_count.imm_val_reg\[10\]
+ _06078_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08745__B1 _03112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ total_design.core.math.pc_val\[3\] total_design.core.program_count.imm_val_reg\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__nor2_1
XANTENNA__08849__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_06730_ total_design.core.regFile.register\[1\]\[4\] net827 net779 total_design.core.regFile.register\[27\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06661_ total_design.core.regFile.register\[15\]\[2\] net604 net581 total_design.core.regFile.register\[6\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a22o_1
XANTENNA__06523__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08400_ total_design.keypad0.key_out\[13\] _03754_ vssd1 vssd1 vccd1 vccd1 _03756_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12057__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06519__D net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09380_ _04617_ _04618_ net701 vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__a21oi_1
X_06592_ total_design.core.regFile.register\[9\]\[1\] net740 net728 net723 vssd1 vssd1
+ vccd1 vccd1 _02163_ sky130_fd_sc_hd__and4_1
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08331_ total_design.core.data_mem.data_write_adr_reg\[23\] net546 net538 total_design.core.data_mem.data_read_adr_reg\[23\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08262_ net1364 net559 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[12\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_117_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07484__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07213_ total_design.core.ctrl.instruction\[25\] net889 vssd1 vssd1 vccd1 vccd1 _02750_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08193_ total_design.core.data_mem.data_write_adr_reg\[29\] total_design.core.data_mem.data_write_adr_reg\[28\]
+ total_design.core.data_mem.data_write_adr_reg\[31\] total_design.core.data_mem.data_write_adr_reg\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__or4_1
XANTENNA__08028__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07236__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07144_ total_design.core.regFile.register\[0\]\[11\] net874 _02671_ _02685_ vssd1
+ vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14471__D net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07075_ total_design.core.regFile.register\[11\]\[10\] net794 net783 total_design.core.regFile.register\[2\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1035_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout495_A _05005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ total_design.core.regFile.register\[3\]\[28\] net867 net820 total_design.core.regFile.register\[17\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10801__B _01852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06762__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ _03598_ net448 net296 _04604_ _04939_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__o221ai_1
X_06928_ total_design.core.regFile.register\[15\]\[7\] net849 net826 total_design.core.regFile.register\[19\]\[7\]
+ _02469_ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__a221o_1
XANTENNA__06279__A net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ _04868_ _04873_ net535 vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06859_ total_design.core.regFile.register\[13\]\[6\] net668 net564 total_design.core.regFile.register\[3\]\[6\]
+ _02401_ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout548_X net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09578_ net705 _04807_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08529_ _03866_ _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11540_ net1794 _05652_ net148 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06218__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11471_ net1566 _05671_ net155 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__mux2_1
XANTENNA__08019__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08941__B _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire458 _02487_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_4
X_10422_ net178 net2158 net386 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__mux2_1
X_13210_ clknet_leaf_132_clk _00677_ net1196 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14190_ clknet_leaf_79_clk _01370_ net1218 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_115_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10353_ net191 net2867 net489 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__mux2_1
X_13141_ clknet_leaf_158_clk _00608_ net1143 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06450__A1 total_design.core.ctrl.instruction\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_143_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13072_ clknet_leaf_185_clk _00539_ net1037 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09519__A2 _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ net201 net1982 net498 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__mux2_1
XANTENNA__06450__B2 total_design.core.ctrl.instruction\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_104_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12023_ total_design.lcd_display.row_1\[89\] _05812_ _05843_ total_design.lcd_display.row_1\[121\]
+ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_163_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08742__A3 _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11095__A _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout580 _02087_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_8
Xfanout591 net592 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10203__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13974_ clknet_leaf_100_clk _01154_ net1237 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_12925_ clknet_leaf_10_clk _00392_ net1019 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12039__B1 _05832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12856_ clknet_leaf_133_clk _00323_ net1195 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06910__C1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11807_ total_design.lcd_display.cnt_20ms\[4\] total_design.lcd_display.cnt_20ms\[5\]
+ _03911_ total_design.lcd_display.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__a31o_1
X_12787_ clknet_leaf_192_clk _00254_ net1032 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14526_ net1298 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
X_11738_ net1653 net957 net290 total_design.core.data_bus_o\[10\] vssd1 vssd1 vccd1
+ vccd1 _01366_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_25_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14457_ clknet_leaf_53_clk net1384 net1095 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09207__A1 _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11669_ _05671_ net1677 net132 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13408_ clknet_leaf_192_clk _00875_ net1032 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07218__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14388_ clknet_leaf_164_clk _01529_ net1164 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08570__C net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13339_ clknet_leaf_144_clk _00806_ net1174 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07900_ total_design.core.regFile.register\[29\]\[26\] net656 net618 total_design.core.regFile.register\[10\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__a22o_1
X_08880_ _04132_ _04133_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09027__X _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07831_ total_design.core.regFile.register\[1\]\[25\] net828 _03332_ _03334_ vssd1
+ vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__a211o_1
XANTENNA__06744__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10113__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07762_ total_design.core.regFile.register\[25\]\[23\] net647 net573 total_design.core.regFile.register\[24\]\[23\]
+ _03258_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09501_ total_design.core.math.pc_val\[20\] _04715_ vssd1 vssd1 vccd1 vccd1 _04735_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09902__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06713_ total_design.core.regFile.register\[7\]\[3\] net651 net604 total_design.core.regFile.register\[15\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__a22o_1
X_07693_ total_design.core.regFile.register\[5\]\[22\] net807 _03189_ _03202_ vssd1
+ vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06644_ net966 _02020_ net888 net967 _02212_ vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[2\]
+ sky130_fd_sc_hd__a221o_2
X_09432_ _04621_ _04668_ net463 vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06575_ net691 _02145_ _02146_ _02147_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__or4_1
X_09363_ net312 _04409_ _04602_ net297 vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__a211o_1
XANTENNA__09446__A1 _02968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06546__B net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08314_ net1502 net940 _03691_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[14\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07457__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ _04193_ _04531_ _04532_ _04533_ _04536_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_23_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_10 total_design.data_in_BUS\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08245_ net1453 net542 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[28\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_74_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout410_A net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1152_A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout129_X net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09349__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08176_ net890 _03090_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[19\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_183_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07127_ total_design.core.regFile.register\[15\]\[11\] net849 net830 total_design.core.regFile.register\[1\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_132_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07058_ total_design.core.regFile.register\[20\]\[10\] net670 net608 total_design.core.regFile.register\[18\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout877_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_198_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06735__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout665_X net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10023__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_121_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09812__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10971_ _05191_ _05197_ _05194_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout832_X net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12710_ clknet_leaf_201_clk _00177_ net1003 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13690_ clknet_leaf_55_clk total_design.core.data_mem.data_read_adr_i\[30\] net1114
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_136_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12641_ clknet_leaf_121_clk _00108_ net1192 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09437__B2 _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07448__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ clknet_leaf_30_clk _00039_ net1064 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11795__A2 _01911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14311_ clknet_leaf_63_clk _01472_ net1124 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_11523_ net1620 _05618_ net145 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10693__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07568__A _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14242_ clknet_leaf_108_clk _01422_ net1228 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11454_ _05674_ _05675_ _05478_ _05480_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__and4b_2
XFILLER_0_135_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10405_ net255 net2468 net385 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__mux2_1
Xwire299 _03177_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__buf_4
X_11385_ net304 net510 _05031_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__or3b_1
X_14173_ clknet_leaf_31_clk _01353_ net1061 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06191__B net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13124_ clknet_leaf_108_clk _00591_ net1223 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10336_ net266 net2619 net491 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11377__X _05636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06974__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10267_ net281 net2049 net496 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__mux2_1
X_13055_ clknet_leaf_183_clk _00522_ net1040 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12006_ total_design.lcd_display.row_1\[40\] _05821_ _05839_ total_design.lcd_display.row_1\[56\]
+ _05867_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__a221o_1
X_10198_ net2873 net392 vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__nand2_1
XANTENNA__09125__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13957_ clknet_leaf_92_clk _01137_ net1262 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07136__C1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11553__A _05478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11483__A1 _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07687__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12908_ clknet_leaf_167_clk _00375_ net1156 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13888_ clknet_leaf_110_clk _01068_ net1227 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12839_ clknet_leaf_18_clk _00306_ net1048 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09428__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07439__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06360_ net951 net950 total_design.core.ctrl.instruction\[23\] net952 vssd1 vssd1
+ vccd1 vccd1 _01936_ sky130_fd_sc_hd__o211a_1
XANTENNA__08862__A total_design.core.instr_fetch vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14509_ net72 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06291_ _01869_ _01861_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08030_ total_design.core.regFile.register\[27\]\[29\] net779 net758 total_design.core.regFile.register\[4\]\[29\]
+ _03513_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__a221o_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire299_X net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold803 total_design.core.regFile.register\[5\]\[16\] vssd1 vssd1 vccd1 vccd1 net2119
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 total_design.core.regFile.register\[27\]\[25\] vssd1 vssd1 vccd1 vccd1 net2130
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10108__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold825 total_design.core.regFile.register\[2\]\[9\] vssd1 vssd1 vccd1 vccd1 net2141
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold836 total_design.core.regFile.register\[9\]\[20\] vssd1 vssd1 vccd1 vccd1 net2152
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold847 total_design.lcd_display.cnt_20ms\[2\] vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07611__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold858 total_design.core.regFile.register\[14\]\[5\] vssd1 vssd1 vccd1 vccd1 net2174
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09981_ net169 net2631 net418 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__mux2_1
Xhold869 total_design.core.regFile.register\[31\]\[20\] vssd1 vssd1 vccd1 vccd1 net2185
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06965__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_75 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08932_ _01746_ _04101_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__nor2_1
X_08863_ _04112_ _04113_ _04116_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__or3_4
Xhold1503 total_design.core.regFile.register\[2\]\[8\] vssd1 vssd1 vccd1 vccd1 net2819
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13716__Q total_design.core.data_cpu_o\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06717__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1514 total_design.core.regFile.register\[0\]\[12\] vssd1 vssd1 vccd1 vccd1 net2830
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1525 total_design.core.regFile.register\[17\]\[12\] vssd1 vssd1 vccd1 vccd1 net2841
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07814_ total_design.core.regFile.register\[12\]\[24\] net567 _03315_ _03318_ vssd1
+ vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__a211o_1
Xhold1536 total_design.core.regFile.register\[21\]\[26\] vssd1 vssd1 vccd1 vccd1 net2852
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1547 total_design.core.regFile.register\[8\]\[20\] vssd1 vssd1 vccd1 vccd1 net2863
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1558 total_design.core.regFile.register\[0\]\[20\] vssd1 vssd1 vccd1 vccd1 net2874
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08794_ total_design.core.data_mem.data_cpu_i\[14\] _02818_ vssd1 vssd1 vccd1 vccd1
+ _04049_ sky130_fd_sc_hd__and2b_1
XFILLER_0_165_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1569 total_design.core.math.pc_val\[13\] vssd1 vssd1 vccd1 vccd1 net2885 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07390__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07941__A total_design.core.data_mem.data_cpu_i\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07745_ total_design.core.regFile.register\[0\]\[23\] net873 _03245_ _03252_ vssd1
+ vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout360_A _05017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06828__Y _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08756__B _03273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11474__A1 _05652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07676_ _03184_ _03186_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__xnor2_4
XANTENNA__07142__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09415_ _04651_ _04652_ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06627_ total_design.core.regFile.register\[1\]\[2\] net830 _02193_ _02196_ vssd1
+ vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout625_A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout246_X net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ net970 net885 net755 total_design.core.data_cpu_o\[13\] vssd1 vssd1 vccd1
+ vccd1 _04587_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06558_ total_design.core.regFile.register\[13\]\[1\] net920 net946 net909 vssd1
+ vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__and4_1
XFILLER_0_164_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08772__A _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ net256 net2249 net453 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06489_ total_design.core.regFile.register\[5\]\[0\] net743 net735 net729 vssd1 vssd1
+ vccd1 vccd1 _02063_ sky130_fd_sc_hd__and4_1
XFILLER_0_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08228_ net1457 net544 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[11\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_62_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07850__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout994_A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08159_ net892 _02241_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[2\]
+ sky130_fd_sc_hd__nor2_1
X_11170_ _05428_ _05415_ _05414_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07602__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09807__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10201__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12969__RESET_B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06956__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ net286 net2002 net398 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10052_ _04118_ _04980_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06231__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06708__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11701__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07381__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13811_ clknet_leaf_71_clk total_design.core.data_mem.data_cpu_i\[20\] net1205 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[20\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10688__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11373__A _05049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11465__A1 _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13742_ clknet_leaf_71_clk total_design.core.data_mem.stored_write_data\[17\] net1206
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[17\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07570__B _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10954_ _05203_ _05197_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07133__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14457__Q total_design.core.instr_mem.instruction_adr_i\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13673_ clknet_leaf_55_clk total_design.core.data_mem.data_read_adr_i\[13\] net1117
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[13\] sky130_fd_sc_hd__dfrtp_1
X_10885_ _05120_ _05125_ _05140_ _05119_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__o22ai_4
Xclkbuf_leaf_191_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_191_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12624_ clknet_leaf_185_clk _00091_ net1037 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12555_ net1449 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06644__A1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11506_ net1829 _05613_ net149 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07841__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12486_ net980 net972 net884 _01697_ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14225_ clknet_leaf_57_clk _01405_ net1115 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dfrtp_1
X_11437_ net1534 _05680_ net159 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14156_ clknet_leaf_31_clk _01336_ net1061 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output87_A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11368_ _05392_ net304 vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__nor2_4
XANTENNA__06947__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13107_ clknet_leaf_180_clk _00574_ net1042 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10319_ net193 net2496 net492 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__mux2_1
X_14087_ clknet_leaf_83_clk _01267_ net1243 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_11299_ _05549_ _05557_ _05550_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__a21o_1
XANTENNA__09346__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13038_ clknet_leaf_190_clk _00505_ net1032 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1150 net1154 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__clkbuf_4
Xfanout1161 net1162 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__clkbuf_2
Xfanout1172 net1265 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__buf_2
Xfanout1183 net1201 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07372__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1194 net1200 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10598__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07530_ total_design.core.regFile.register\[25\]\[19\] net648 net602 total_design.core.regFile.register\[31\]\[19\]
+ _03046_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07124__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07461_ total_design.core.regFile.register\[16\]\[17\] _01932_ net831 total_design.core.regFile.register\[31\]\[17\]
+ net691 vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_182_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_182_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_83_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09200_ _04431_ _04445_ _04446_ net451 vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__a31o_1
X_06412_ net926 net914 net912 vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07392_ total_design.core.regFile.register\[4\]\[16\] net815 net808 total_design.core.regFile.register\[5\]\[16\]
+ net693 vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09040__X _04292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11759__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09131_ net322 _04243_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__nor2_1
X_06343_ net971 net973 total_design.core.ctrl.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ _01919_ sky130_fd_sc_hd__and3b_1
XFILLER_0_151_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08085__B1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09282__C1 _04105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09062_ total_design.core.data_cpu_o\[2\] net757 net905 total_design.core.math.pc_val\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__o2bb2a_1
X_06274_ total_design.core.instr_mem.instruction_adr_i\[2\] total_design.core.instr_mem.instruction_adr_stored\[2\]
+ net984 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08013_ _03416_ _03420_ _03463_ _03464_ _03509_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__o311a_1
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09034__C1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold600 total_design.core.regFile.register\[16\]\[22\] vssd1 vssd1 vccd1 vccd1 net1916
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout206_A _04740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold611 total_design.core.regFile.register\[9\]\[30\] vssd1 vssd1 vccd1 vccd1 net1927
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 total_design.core.regFile.register\[20\]\[20\] vssd1 vssd1 vccd1 vccd1 net1938
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 total_design.core.regFile.register\[21\]\[25\] vssd1 vssd1 vccd1 vccd1 net1949
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 total_design.core.regFile.register\[31\]\[23\] vssd1 vssd1 vccd1 vccd1 net1960
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06840__A total_design.core.ctrl.instruction\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold655 total_design.core.regFile.register\[24\]\[27\] vssd1 vssd1 vccd1 vccd1 net1971
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10195__A1 _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07596__C1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold666 total_design.core.regFile.register\[14\]\[21\] vssd1 vssd1 vccd1 vccd1 net1982
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold677 total_design.core.regFile.register\[9\]\[28\] vssd1 vssd1 vccd1 vccd1 net1993
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold688 total_design.core.regFile.register\[2\]\[12\] vssd1 vssd1 vccd1 vccd1 net2004
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 total_design.keypad0.counter\[14\] vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09964_ net236 net2029 net421 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__mux2_1
X_08915_ net471 _03322_ _04168_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__o21bai_1
X_09895_ net242 net2738 net429 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout575_A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1300 total_design.core.regFile.register\[1\]\[5\] vssd1 vssd1 vccd1 vccd1 net2616
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1311 total_design.core.regFile.register\[24\]\[10\] vssd1 vssd1 vccd1 vccd1 net2627
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 total_design.core.regFile.register\[29\]\[31\] vssd1 vssd1 vccd1 vccd1 net2638
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07899__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ total_design.core.ctrl.instruction\[12\] _01747_ _02029_ vssd1 vssd1 vccd1
+ vccd1 _04101_ sky130_fd_sc_hd__or3b_2
Xhold1333 total_design.keypad0.counter\[12\] vssd1 vssd1 vccd1 vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1344 total_design.core.regFile.register\[0\]\[7\] vssd1 vssd1 vccd1 vccd1 net2660
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1355 total_design.data_in_BUS\[3\] vssd1 vssd1 vccd1 vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 total_design.core.regFile.register\[13\]\[17\] vssd1 vssd1 vccd1 vccd1 net2682
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1377 total_design.core.regFile.register\[17\]\[25\] vssd1 vssd1 vccd1 vccd1 net2693
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout742_A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ _04022_ _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__nand2_1
XANTENNA__06571__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1388 total_design.core.data_bus_o\[1\] vssd1 vssd1 vccd1 vccd1 net2704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1399 total_design.core.regFile.register\[11\]\[0\] vssd1 vssd1 vccd1 vccd1 net2715
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11447__A1 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07728_ total_design.core.regFile.register\[17\]\[23\] net819 net779 total_design.core.regFile.register\[27\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__a22o_1
XANTENNA__10301__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06287__A net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07115__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11998__A2 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07659_ total_design.core.regFile.register\[16\]\[21\] net634 net605 total_design.core.regFile.register\[15\]\[21\]
+ _03169_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_173_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_173_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_101_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10670_ net240 net2683 net361 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09329_ net701 _04569_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_11_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12340_ total_design.core.math.pc_val\[22\] total_design.core.program_count.imm_val_reg\[22\]
+ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout997_X net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12271_ net895 _06111_ net524 vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ clknet_leaf_84_clk _01190_ net1249 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_79_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11222_ _05372_ _05378_ _05362_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a21boi_1
XANTENNA__06929__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11153_ _05411_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__inv_2
X_10104_ net213 net2779 net402 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__mux2_1
XANTENNA__11087__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11084_ net351 _05280_ _05290_ _05292_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10035_ net224 net2212 net412 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__mux2_1
XANTENNA__08000__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07354__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11438__A1 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10211__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11986_ net474 _05842_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__nor2_4
XFILLER_0_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07106__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13725_ clknet_leaf_114_clk total_design.core.data_mem.stored_write_data\[0\] net1207
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[0\] sky130_fd_sc_hd__dfrtp_1
X_10937_ _05161_ _05192_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_164_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_164_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13656_ clknet_leaf_56_clk total_design.core.data_mem.data_write_adr_i\[28\] net1113
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10868_ _05107_ _05126_ _05121_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12607_ clknet_leaf_183_clk _00074_ net1136 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08067__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ clknet_leaf_32_clk total_design.core.data_mem.data_bus_i\[23\] net1063 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[23\] sky130_fd_sc_hd__dfrtp_1
X_10799_ total_design.core.data_bus_o\[13\] _05028_ vssd1 vssd1 vccd1 vccd1 _05058_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12538_ total_design.core.ctrl.instruction\[31\] net885 _02149_ _03091_ net550 vssd1
+ vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[22\] sky130_fd_sc_hd__a221o_1
XFILLER_0_81_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06363__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12469_ net2305 _01686_ _01688_ _01689_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__o211a_1
X_14208_ clknet_leaf_60_clk _01388_ net1131 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12166__A2 _02241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14139_ clknet_leaf_89_clk _01319_ net1260 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout409 _04987_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07593__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ total_design.core.regFile.register\[28\]\[8\] net587 _02509_ _02511_ vssd1
+ vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__a211o_1
X_08700_ _03954_ _03967_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09680_ total_design.core.math.pc_val\[27\] _04861_ total_design.core.math.pc_val\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_33_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06892_ total_design.core.ctrl.instruction\[19\] net885 vssd1 vssd1 vccd1 vccd1 _02447_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07345__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08631_ total_design.lcd_display.cnt_500hz\[1\] total_design.lcd_display.cnt_500hz\[0\]
+ total_design.lcd_display.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_85_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10121__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08562_ net1847 net338 net718 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[17\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__09910__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13797__CLK clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07513_ _03029_ _03030_ _03032_ _03033_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08493_ _03713_ _03771_ _03844_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_155_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_155_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout156_A _05681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07444_ total_design.core.regFile.register\[0\]\[17\] net682 _02962_ _02967_ vssd1
+ vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__o22a_4
XFILLER_0_174_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07375_ _02900_ _02901_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1065_A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09114_ _04146_ _04151_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__and2b_1
X_06326_ net512 _01904_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__and2_1
XANTENNA__07805__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06257_ total_design.core.data_adr_o\[11\] _01835_ net963 vssd1 vssd1 vccd1 vccd1
+ _01836_ sky130_fd_sc_hd__mux2_1
X_09045_ _04296_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1232_A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06188_ _01725_ net1266 net1087 total_design.core.mem_ctrl.state\[2\] total_design.core.mem_ctrl.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__a311o_1
Xhold430 total_design.lcd_display.row_2\[94\] vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 total_design.lcd_display.row_2\[40\] vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold452 total_design.lcd_display.row_2\[92\] vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout692_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold463 total_design.lcd_display.row_2\[24\] vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13818__D total_design.core.data_mem.data_cpu_i\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 net57 vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 total_design.lcd_display.row_1\[124\] vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold496 net59 vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07584__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout910 _01950_ vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout921 net924 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__buf_1
XFILLER_0_99_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout932 total_design.keypad0.key_out\[12\] vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__buf_2
XFILLER_0_25_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09947_ net171 net2450 net422 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__mux2_1
Xfanout943 _03674_ vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout480_X net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout954 net955 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__buf_2
XANTENNA__06792__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout957_A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_X net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_146_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout965 total_design.core.ctrl.instruction\[23\] vssd1 vssd1 vccd1 vccd1 net965
+ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout976 net978 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__buf_2
XANTENNA__10820__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout987 total_design.keypad0.key_clk vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__clkbuf_2
X_09878_ net175 net2095 net431 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__mux2_1
Xfanout998 total_design.core.data_mem.data_read vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 total_design.core.regFile.register\[15\]\[25\] vssd1 vssd1 vccd1 vccd1 net2446
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 total_design.core.regFile.register\[14\]\[20\] vssd1 vssd1 vccd1 vccd1 net2457
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07336__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09730__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1152 total_design.core.regFile.register\[10\]\[10\] vssd1 vssd1 vccd1 vccd1 net2468
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ _04036_ _04049_ _04083_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__or3_1
Xhold1163 total_design.core.regFile.register\[16\]\[24\] vssd1 vssd1 vccd1 vccd1 net2479
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1174 total_design.core.regFile.register\[29\]\[4\] vssd1 vssd1 vccd1 vccd1 net2490
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 total_design.core.regFile.register\[23\]\[5\] vssd1 vssd1 vccd1 vccd1 net2501
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 total_design.core.regFile.register\[25\]\[22\] vssd1 vssd1 vccd1 vccd1 net2512
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ total_design.lcd_display.currentState\[4\] total_design.lcd_display.currentState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__nand2_1
XANTENNA__10031__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09820__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12093__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ net1559 net956 _05700_ _01865_ vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_146_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_146_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ clknet_leaf_199_clk _00977_ net1007 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10722_ net166 net1995 net360 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14490_ clknet_leaf_33_clk _01557_ net1070 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_172_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08049__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13441_ clknet_leaf_120_clk _00908_ net1170 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10653_ net178 net2115 net477 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13372_ clknet_leaf_30_clk _00839_ net1064 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10584_ net192 net2399 net371 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__mux2_1
Xclkload19 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_90_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12323_ _01588_ _01589_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12148__A2 _05829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12254_ net897 _06096_ net527 vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11205_ _05442_ _05446_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12185_ net902 _02395_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10206__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11136_ _05390_ _05393_ _05394_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_79_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11108__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ net350 _05280_ _05285_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__or3b_1
XANTENNA__07327__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _04968_ _04980_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11969_ _05746_ _05749_ _05811_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__or3_2
Xclkbuf_leaf_137_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_137_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_169_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_88_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13708_ clknet_leaf_27_clk total_design.core.data_mem.stored_read_data\[15\] net1075
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08573__C net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07103__X _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13639_ clknet_leaf_67_clk total_design.core.data_mem.data_write_adr_i\[11\] net1111
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07160_ total_design.core.ctrl.instruction\[24\] net889 _02698_ net550 vssd1 vssd1
+ vccd1 vccd1 total_design.core.ctrl.imm_32\[12\] sky130_fd_sc_hd__a211o_1
XFILLER_0_26_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11595__A0 _05663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07091_ _02613_ _02633_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06471__C1 total_design.core.ctrl.instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__06390__A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10116__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout206 _04740_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_1
Xfanout217 _04699_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_1
X_09801_ net205 net2592 net438 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__mux2_1
XANTENNA__09905__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout228 net231 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_2
X_07993_ total_design.core.regFile.register\[7\]\[28\] net653 net634 total_design.core.regFile.register\[16\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__a22o_1
Xfanout239 _04564_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_52_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09732_ net467 _04263_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__nand2_1
X_06944_ total_design.core.ctrl.instruction\[20\] net889 _02028_ total_design.core.ctrl.instruction\[28\]
+ _02495_ vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[8\] sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_2_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09663_ _04121_ _04889_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__nor2_1
X_06875_ total_design.core.regFile.register\[15\]\[6\] net848 net769 total_design.core.regFile.register\[7\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a22o_1
X_08614_ net113 net112 net114 net115 vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__and4b_1
X_09594_ _03303_ _03322_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09640__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08545_ _03768_ _03892_ _03893_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout440_A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_128_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1182_A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout159_X net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_A _03676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ total_design.keypad0.key_out\[10\] _03828_ vssd1 vssd1 vccd1 vccd1 _03829_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__08109__X _03602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07427_ total_design.core.regFile.register\[6\]\[17\] net581 net577 total_design.core.regFile.register\[27\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout705_A _04204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07358_ _02877_ _02881_ _02887_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06309_ _01872_ _01887_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__nor2_4
XANTENNA__07667__Y _03178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07254__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07289_ total_design.core.regFile.register\[8\]\[14\] net802 _01986_ total_design.core.regFile.register\[2\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09028_ net506 _04280_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__and2_1
XANTENNA__06462__C1 total_design.core.ctrl.instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_20_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold260 total_design.lcd_display.row_1\[51\] vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10026__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold271 net92 vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 total_design.lcd_display.row_1\[42\] vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07557__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold293 net81 vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout862_X net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06765__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout740 net743 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__clkbuf_2
Xfanout751 net752 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__clkbuf_4
Xfanout762 _01999_ vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__buf_4
X_13990_ clknet_leaf_96_clk _01170_ net1254 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout773 net774 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__buf_4
Xfanout784 net785 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__buf_4
Xfanout795 net797 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09703__B1 _04924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ clknet_leaf_0_clk _00408_ net1003 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_161_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12872_ clknet_leaf_117_clk _00339_ net1159 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07190__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11823_ net1870 _05713_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__xor2_1
XANTENNA__10696__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_119_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14542_ net1314 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_0_68_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11754_ net91 net960 net293 total_design.core.data_bus_o\[26\] vssd1 vssd1 vccd1
+ vccd1 _01382_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10705_ net229 net2639 net358 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__mux2_1
X_14473_ clknet_leaf_38_clk _01540_ net1079 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11685_ wishbone.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__and2_1
X_13424_ clknet_leaf_190_clk _00891_ net1034 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10636_ net253 net2669 net476 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__mux2_1
XANTENNA__11577__A0 _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload108 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 clkload108/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload119 clknet_leaf_169_clk vssd1 vssd1 vccd1 vccd1 clkload119/Y sky130_fd_sc_hd__inv_6
XFILLER_0_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13355_ clknet_leaf_107_clk _00822_ net1224 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10567_ net267 net1957 net370 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12306_ _06132_ _01574_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__or2_1
XANTENNA__07796__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08993__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13286_ clknet_leaf_199_clk _00753_ net1001 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10498_ net283 net2293 net480 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__mux2_1
X_12237_ total_design.core.math.pc_val\[10\] net527 _06075_ _06081_ vssd1 vssd1 vccd1
+ vccd1 _01480_ sky130_fd_sc_hd__a22o_1
XANTENNA__07548__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08745__A1 _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08745__B2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12168_ total_design.core.math.pc_val\[3\] total_design.core.program_count.imm_val_reg\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__and2_1
XANTENNA__06756__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11119_ _05376_ _05377_ _05371_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__a21oi_4
X_12099_ total_design.lcd_display.row_1\[85\] _05815_ _05838_ total_design.lcd_display.row_1\[29\]
+ _05955_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06369__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06660_ total_design.core.regFile.register\[7\]\[2\] net651 _02227_ net686 vssd1
+ vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a211o_1
XANTENNA__07181__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06591_ total_design.core.regFile.register\[28\]\[1\] net744 net738 net726 vssd1
+ vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__and4_1
XFILLER_0_143_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10068__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08330_ net1470 net938 _03699_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[22\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08261_ net1363 net559 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[11\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_89_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07212_ _02747_ _02748_ net722 vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__a21oi_1
X_08192_ total_design.core.data_mem.data_write_adr_reg\[25\] total_design.core.data_mem.data_write_adr_reg\[24\]
+ total_design.core.data_mem.data_write_adr_reg\[27\] total_design.core.data_mem.data_write_adr_reg\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__or4_1
XANTENNA__11568__A0 _05655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07143_ _02673_ _02675_ _02677_ _02684_ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__or4_1
XFILLER_0_160_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06832__B _02367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07787__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07074_ total_design.core.regFile.register\[8\]\[10\] net802 net767 total_design.core.regFile.register\[7\]\[10\]
+ _02618_ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__a221o_1
XANTENNA__13719__Q total_design.core.data_cpu_o\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08105__A _03595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06551__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07539__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout390_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11740__B1 _05049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ total_design.core.regFile.register\[29\]\[28\] net799 _03470_ _03473_ vssd1
+ vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__a211o_1
X_09715_ net969 _03598_ _03599_ _04100_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__o211ai_1
X_06927_ total_design.core.regFile.register\[26\]\[7\] net872 net813 total_design.core.regFile.register\[23\]\[7\]
+ _02480_ vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout655_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ net704 _04870_ _04871_ _04872_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__or4b_1
X_06858_ total_design.core.regFile.register\[20\]\[6\] net672 net606 total_design.core.regFile.register\[15\]\[6\]
+ _02400_ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__a221o_1
XANTENNA__07172__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07711__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09577_ _03277_ _04762_ _04785_ _03326_ _03275_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__o311a_1
XANTENNA__09449__C1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06789_ total_design.core.regFile.register\[9\]\[5\] net665 net634 total_design.core.regFile.register\[16\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08528_ _03861_ _03877_ _03876_ _03875_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_33_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07475__A1 total_design.core.ctrl.instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08459_ _03777_ _03783_ _03812_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout610_X net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11470_ net1751 _05680_ net156 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_6__f_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14411__RESET_B net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11559__A0 _05626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10421_ net182 net2799 net387 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__mux2_1
XANTENNA__12220__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10231__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07778__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13140_ clknet_leaf_143_clk _00607_ net1175 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10352_ net193 net2336 net488 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10782__A1 total_design.core.data_bus_o\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06461__C net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13071_ clknet_leaf_147_clk _00538_ net1152 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10283_ net208 net2457 net496 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__mux2_1
X_12022_ total_design.lcd_display.row_2\[65\] _05819_ _05849_ total_design.lcd_display.row_2\[49\]
+ _05882_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_163_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06738__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout570 _02091_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07950__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout581 _02085_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_8
Xfanout592 _02081_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__buf_4
X_13973_ clknet_leaf_91_clk _01153_ net1262 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09152__A1 total_design.core.data_cpu_o\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ clknet_leaf_30_clk _00391_ net1060 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07163__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07702__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12855_ clknet_leaf_166_clk _00322_ net1157 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11806_ total_design.lcd_display.cnt_20ms\[4\] total_design.lcd_display.cnt_20ms\[5\]
+ total_design.lcd_display.cnt_20ms\[6\] _03911_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__and4_1
XFILLER_0_139_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12786_ clknet_leaf_137_clk _00253_ net1179 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08112__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11798__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14195__Q net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14525_ net1297 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XANTENNA__07466__A1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11737_ net1840 net957 _05077_ _05695_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14456_ clknet_leaf_53_clk net1485 net1109 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11668_ _05680_ net1721 net131 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__mux2_1
XANTENNA__09207__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13407_ clknet_leaf_184_clk _00874_ net1039 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12211__A1 _02016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08415__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10619_ net182 net2317 net366 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__mux2_1
X_14387_ clknet_leaf_152_clk _01528_ net1139 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11599_ _05632_ net1582 net139 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10222__A0 _04909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13338_ clknet_leaf_125_clk _00805_ net1190 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06977__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06371__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13269_ clknet_leaf_157_clk _00736_ net1140 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12514__A2 total_design.core.ctrl.instruction\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08212__X _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06729__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ total_design.core.regFile.register\[30\]\[25\] net839 net768 total_design.core.regFile.register\[7\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__a22o_1
X_07761_ total_design.core.regFile.register\[15\]\[23\] net604 _03267_ net686 vssd1
+ vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09500_ net449 _04733_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__nor2_1
X_06712_ total_design.core.regFile.register\[2\]\[3\] net637 net621 total_design.core.regFile.register\[4\]\[3\]
+ _02276_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__a221o_1
X_07692_ total_design.core.regFile.register\[20\]\[22\] net816 net799 total_design.core.regFile.register\[29\]\[22\]
+ _03188_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09431_ _04218_ _04256_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__nand2_1
X_06643_ total_design.core.ctrl.instruction\[9\] _01918_ _02149_ _01738_ vssd1 vssd1
+ vccd1 vccd1 _02212_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06901__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09362_ net312 _04412_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__nor2_1
X_06574_ total_design.core.regFile.register\[3\]\[1\] net865 net853 total_design.core.regFile.register\[28\]\[1\]
+ _02123_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a221o_1
XANTENNA__11789__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08313_ total_design.core.data_mem.data_write_adr_reg\[14\] net548 net540 total_design.core.data_mem.data_read_adr_reg\[14\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09293_ _02693_ net508 net298 _04534_ _04535_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__o221ai_4
XANTENNA_11 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout236_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08244_ net1483 net542 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[27\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_43_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11687__A_N total_design.bus_full vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08175_ net890 _03040_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[18\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06680__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout403_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10213__A0 _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06562__B net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07126_ total_design.core.regFile.register\[14\]\[11\] net861 net764 total_design.core.regFile.register\[6\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_132_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07057_ total_design.core.regFile.register\[30\]\[10\] net659 _02601_ vssd1 vssd1
+ vccd1 vccd1 _02602_ sky130_fd_sc_hd__a21o_1
XANTENNA__06432__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09906__A0 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_A _01995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10304__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__B1 _01995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ _03443_ _03446_ _03456_ _03457_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ _05191_ _05194_ _05197_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__or3_1
XANTENNA_hold448_A total_design.core.math.pc_val\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09629_ _03418_ net509 _04687_ _04693_ _04856_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_67_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ clknet_leaf_191_clk _00107_ net1032 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12571_ net1412 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_156_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_50_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14310_ clknet_leaf_103_clk _00010_ net1238 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11522_ net1833 _05621_ net145 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07999__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14241_ clknet_leaf_108_clk _01421_ net1228 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11453_ net1585 _05630_ net159 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__mux2_1
XANTENNA__06472__B net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10204__A0 _04563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ net249 net2769 net387 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__mux2_1
X_14172_ clknet_leaf_32_clk _01352_ net1066 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11384_ _05586_ _05642_ _05640_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__o21a_2
XFILLER_0_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06959__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13123_ clknet_leaf_9_clk _00590_ net1019 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10335_ net274 net2843 net490 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13054_ clknet_leaf_180_clk _00521_ net1044 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10266_ net268 net2831 net496 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__mux2_1
X_12005_ total_design.lcd_display.row_1\[80\] _05815_ _05830_ total_design.lcd_display.row_1\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09373__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10197_ _04451_ net390 _04995_ vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07384__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07923__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11393__X _05652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13956_ clknet_leaf_98_clk _01136_ net1244 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07136__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06487__X _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11553__B _05479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12907_ clknet_leaf_108_clk _00374_ net1224 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13887_ clknet_leaf_82_clk _01067_ net1220 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12838_ clknet_leaf_199_clk _00305_ net1001 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12769_ clknet_leaf_121_clk _00236_ net1170 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08100__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14508_ net72 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
X_06290_ _01866_ _01868_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14439_ clknet_leaf_59_clk net1560 net1127 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06662__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06382__B net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09061__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold804 total_design.core.regFile.register\[9\]\[23\] vssd1 vssd1 vccd1 vccd1 net2120
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 total_design.core.regFile.register\[29\]\[11\] vssd1 vssd1 vccd1 vccd1 net2131
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 total_design.core.regFile.register\[26\]\[26\] vssd1 vssd1 vccd1 vccd1 net2142
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold837 total_design.core.regFile.register\[28\]\[29\] vssd1 vssd1 vccd1 vccd1 net2153
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold848 total_design.core.regFile.register\[18\]\[20\] vssd1 vssd1 vccd1 vccd1 net2164
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09980_ net172 net2811 net420 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold859 total_design.core.regFile.register\[15\]\[5\] vssd1 vssd1 vccd1 vccd1 net2175
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08931_ net508 net533 _02118_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10124__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08862_ total_design.core.instr_fetch _04114_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__or2_2
Xhold1504 total_design.core.regFile.register\[27\]\[14\] vssd1 vssd1 vccd1 vccd1 net2820
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1515 total_design.core.regFile.register\[14\]\[3\] vssd1 vssd1 vccd1 vccd1 net2831
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07813_ total_design.core.regFile.register\[8\]\[24\] net594 _03316_ _03317_ vssd1
+ vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__a211o_1
Xhold1526 total_design.core.regFile.register\[22\]\[21\] vssd1 vssd1 vccd1 vccd1 net2842
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09913__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1537 total_design.core.regFile.register\[19\]\[0\] vssd1 vssd1 vccd1 vccd1 net2853
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08793_ total_design.core.data_mem.data_cpu_i\[12\] _02718_ vssd1 vssd1 vccd1 vccd1
+ _04048_ sky130_fd_sc_hd__and2b_1
XFILLER_0_93_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1548 total_design.lcd_display.cnt_500hz\[7\] vssd1 vssd1 vccd1 vccd1 net2864
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1559 total_design.core.regFile.register\[0\]\[25\] vssd1 vssd1 vccd1 vccd1 net2875
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07744_ _03247_ _03248_ _03249_ _03251_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_88_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07127__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12120__B1 _05839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13732__Q total_design.core.data_bus_o\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ _03093_ _03136_ _03134_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout353_A _05018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06557__B net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09414_ total_design.core.math.pc_val\[15\] _04609_ total_design.core.math.pc_val\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_45_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06626_ total_design.core.regFile.register\[17\]\[2\] net819 _02194_ _02195_ vssd1
+ vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ net904 _04585_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout520_A _01885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06557_ total_design.core.regFile.register\[23\]\[1\] net925 net911 net907 vssd1
+ vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout141_X net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout239_X net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08772__B _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09220__Y _04466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09276_ _04515_ _04519_ net452 vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__a21oi_4
X_06488_ net740 net735 net728 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_134_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08227_ net1393 net543 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[10\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__06653__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08158_ net892 _02188_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[1\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_151_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07063__C1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07109_ total_design.core.regFile.register\[9\]\[11\] _02049_ net633 total_design.core.regFile.register\[16\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08089_ total_design.core.regFile.register\[20\]\[30\] net672 net591 total_design.core.regFile.register\[1\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10120_ _04115_ _04989_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__nand2_4
XFILLER_0_101_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_99_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_42_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09355__A1 _02845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ net163 net2086 net411 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__mux2_1
XANTENNA__10034__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07905__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09823__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ clknet_leaf_113_clk total_design.core.data_mem.data_cpu_i\[19\] net1206 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[19\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07118__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12111__B1 _05912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08315__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13741_ clknet_leaf_72_clk total_design.core.data_mem.stored_write_data\[16\] net1205
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10953_ _05211_ _05200_ _05178_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06467__B net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13672_ clknet_leaf_58_clk total_design.core.data_mem.data_read_adr_i\[12\] net1120
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10884_ _05132_ _05138_ _05140_ _05141_ _05129_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_85_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12623_ clknet_leaf_146_clk _00090_ net1178 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_14_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12554_ net1432 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_14_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13797__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11505_ net1533 _05657_ net150 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__mux2_1
X_12485_ net979 net2732 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__and2b_1
XANTENNA__10209__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14224_ clknet_leaf_57_clk _01404_ net1116 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07866__X _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11436_ _05459_ _05629_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__and2_2
XFILLER_0_110_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14155_ clknet_leaf_34_clk _01335_ net1066 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11367_ _05411_ net303 _05625_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__o21a_2
XFILLER_0_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ clknet_leaf_138_clk _00573_ net1184 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_60_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10318_ net197 net2418 net493 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__mux2_1
X_14086_ clknet_leaf_101_clk _01266_ net1237 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_11298_ net248 _05543_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09346__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08149__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13037_ clknet_leaf_4_clk _00504_ net1023 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10249_ net211 net2461 net501 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__mux2_1
XANTENNA__09018__B _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1140 net1141 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__clkbuf_4
Xfanout1151 net1154 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__buf_2
Xfanout1162 net1163 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__clkbuf_2
Xfanout1173 net1181 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__clkbuf_4
Xfanout1184 net1185 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08857__B _02014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1195 net1200 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_117_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07109__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12102__B1 _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_182_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06580__A1 total_design.core.ctrl.instruction\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__06580__B2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08576__C net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13939_ clknet_leaf_93_clk _01119_ net1255 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_62_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07460_ total_design.core.regFile.register\[18\]\[17\] net857 net850 total_design.core.regFile.register\[9\]\[17\]
+ _02973_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08873__A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09321__X _04563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06411_ total_design.core.regFile.register\[2\]\[0\] net923 net948 net917 vssd1 vssd1
+ vccd1 vccd1 _01987_ sky130_fd_sc_hd__and4_1
XANTENNA__12405__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_197_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07391_ _02917_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__inv_2
XANTENNA__11503__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_14_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09130_ _02395_ net705 _04378_ net535 vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__a211o_1
X_06342_ _01915_ _01917_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_40_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09061_ _04292_ _04312_ net451 vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06273_ _01806_ _01818_ _01834_ _01851_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__nand4_4
XANTENNA__06635__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08012_ _03507_ _03508_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__nor2_1
XANTENNA__09908__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold601 total_design.core.regFile.register\[11\]\[27\] vssd1 vssd1 vccd1 vccd1 net1917
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold612 total_design.lcd_display.row_2\[82\] vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold623 total_design.core.regFile.register\[6\]\[7\] vssd1 vssd1 vccd1 vccd1 net1939
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 total_design.core.regFile.register\[10\]\[13\] vssd1 vssd1 vccd1 vccd1 net1950
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 total_design.core.regFile.register\[23\]\[14\] vssd1 vssd1 vccd1 vccd1 net1961
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 total_design.core.regFile.register\[10\]\[21\] vssd1 vssd1 vccd1 vccd1 net1972
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10195__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11392__B2 _05037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold667 total_design.core.regFile.register\[3\]\[1\] vssd1 vssd1 vccd1 vccd1 net1983
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold678 total_design.core.regFile.register\[10\]\[22\] vssd1 vssd1 vccd1 vccd1 net1994
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07060__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09963_ net240 net2191 net418 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_135_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold689 total_design.core.regFile.register\[6\]\[9\] vssd1 vssd1 vccd1 vccd1 net2005
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ net335 _03369_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1010_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ net255 net2177 net426 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__mux2_1
XANTENNA__07348__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1108_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1301 total_design.core.regFile.register\[12\]\[25\] vssd1 vssd1 vccd1 vccd1 net2617
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1312 total_design.core.regFile.register\[25\]\[30\] vssd1 vssd1 vccd1 vccd1 net2628
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08845_ total_design.core.ctrl.instruction\[12\] net967 _02029_ vssd1 vssd1 vccd1
+ vccd1 _04100_ sky130_fd_sc_hd__and3b_2
XANTENNA__11695__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1323 total_design.core.regFile.register\[1\]\[13\] vssd1 vssd1 vccd1 vccd1 net2639
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1334 total_design.core.regFile.register\[22\]\[30\] vssd1 vssd1 vccd1 vccd1 net2650
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout470_A _02111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1345 total_design.core.regFile.register\[13\]\[2\] vssd1 vssd1 vccd1 vccd1 net2661
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout568_A _02092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1356 total_design.core.regFile.register\[16\]\[17\] vssd1 vssd1 vccd1 vccd1 net2672
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1367 total_design.core.regFile.register\[2\]\[11\] vssd1 vssd1 vccd1 vccd1 net2683
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08776_ _04029_ _04030_ _04026_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__and3b_1
Xhold1378 total_design.core.regFile.register\[18\]\[29\] vssd1 vssd1 vccd1 vccd1 net2694
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_108_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1389 _01357_ vssd1 vssd1 vccd1 vccd1 net2705 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07016__X _02564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__B _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07727_ total_design.core.regFile.register\[20\]\[23\] net818 net810 total_design.core.regFile.register\[23\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08312__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07658_ total_design.core.regFile.register\[14\]\[21\] net625 net583 total_design.core.regFile.register\[6\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08783__A _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06609_ total_design.core.regFile.register\[6\]\[1\] net582 _02179_ net689 vssd1
+ vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_101_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06874__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout902_A _02016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07589_ total_design.core.regFile.register\[21\]\[20\] net597 net589 total_design.core.regFile.register\[1\]\[20\]
+ _03102_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1265_X net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10818__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09328_ _04565_ _04566_ _04568_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_153_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14293__Q net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06626__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ _04136_ _04139_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10029__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_117_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09818__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ net993 _04611_ _06109_ _06110_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout892_X net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ _05479_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07587__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ net513 _05154_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__nand2_2
XANTENNA__07051__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10103_ net221 net2615 net403 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11083_ _05285_ _05290_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__nand2_1
XANTENNA__07339__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ net233 net2484 net413 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__mux2_1
XANTENNA__10699__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11985_ net531 _05836_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__nor2_4
XANTENNA__08303__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10936_ _05183_ _05188_ _05190_ _05192_ _05193_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__a2111o_1
X_13724_ clknet_leaf_27_clk total_design.core.data_mem.stored_read_data\[31\] net1077
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[31\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07511__B1 _01992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13655_ clknet_leaf_50_clk total_design.core.data_mem.data_write_adr_i\[27\] net1100
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[27\] sky130_fd_sc_hd__dfrtp_1
X_10867_ _05118_ _05119_ _05125_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06865__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12606_ clknet_leaf_173_clk _00073_ net1056 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08843__D _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13586_ clknet_leaf_33_clk total_design.core.data_mem.data_bus_i\[22\] net1063 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[22\] sky130_fd_sc_hd__dfrtp_1
X_10798_ net350 _05055_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__or2_2
XFILLER_0_82_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12537_ _01730_ net1476 _01888_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12468_ total_design.keypad0.next_rows\[1\] _03983_ _05783_ _03984_ vssd1 vssd1 vccd1
+ vccd1 _01689_ sky130_fd_sc_hd__o31a_1
XFILLER_0_124_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07290__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06941__A total_design.core.ctrl.instruction\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_2_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11419_ net1854 _05344_ _05354_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__mux2_1
X_14207_ clknet_leaf_111_clk _01387_ net1208 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_2
X_12399_ _01656_ _01657_ vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__nand2_1
XANTENNA__11374__A1 total_design.core.data_bus_o\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14138_ clknet_leaf_87_clk _01318_ net1248 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14069_ clknet_leaf_91_clk _01249_ net1263 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[87\]
+ sky130_fd_sc_hd__dfrtp_1
X_06960_ total_design.core.regFile.register\[30\]\[8\] net661 _02497_ _02510_ vssd1
+ vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_3_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06891_ _02312_ _02445_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_33_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08630_ total_design.lcd_display.cnt_500hz\[1\] total_design.lcd_display.cnt_500hz\[0\]
+ total_design.lcd_display.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__a21o_1
XANTENNA__10402__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07750__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08561_ total_design.data_in_BUS\[16\] net340 net719 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[16\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_89_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07512_ total_design.core.regFile.register\[16\]\[18\] net854 _03019_ net691 vssd1
+ vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_18_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08492_ total_design.keypad0.key_out\[13\] net931 total_design.keypad0.key_out\[15\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__or4_1
XANTENNA__07502__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07443_ _02953_ _02964_ _02965_ _02966_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__or4_1
XANTENNA__06856__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout149_A _05682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07374_ total_design.core.regFile.register\[30\]\[16\] net661 net572 total_design.core.regFile.register\[17\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06554__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09113_ net460 _04287_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__nor2_1
X_06325_ _01872_ _01903_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__or2_4
XFILLER_0_127_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06608__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1058_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09044_ _04293_ _04295_ net330 vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__mux2_2
X_06256_ total_design.core.instr_mem.instruction_adr_i\[11\] total_design.core.instr_mem.instruction_adr_stored\[11\]
+ net983 vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__mux2_1
XANTENNA__07281__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09558__A1 _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold420 total_design.lcd_display.row_2\[99\] vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 total_design.lcd_display.row_2\[20\] vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
X_06187_ net998 total_design.core.instr_fetch vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold442 total_design.lcd_display.row_2\[18\] vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 total_design.lcd_display.row_2\[73\] vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold464 total_design.lcd_display.row_2\[36\] vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07033__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold475 total_design.lcd_display.row_2\[44\] vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold486 total_design.lcd_display.row_1\[126\] vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11619__D _05675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout900 net901 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout685_A _02035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold497 total_design.lcd_display.row_2\[126\] vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 net912 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout922 net923 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__clkbuf_2
X_09946_ net174 net2334 net423 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout933 total_design.keypad0.key_out\[9\] vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__buf_2
XFILLER_0_99_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout944 _03674_ vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_4
Xfanout955 _01911_ vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_2
Xfanout966 total_design.core.ctrl.instruction\[22\] vssd1 vssd1 vccd1 vccd1 net966
+ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout977 net978 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1120 total_design.core.regFile.register\[8\]\[7\] vssd1 vssd1 vccd1 vccd1 net2436
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09877_ net178 net2266 net432 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout852_A _01951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout988 total_design.core.program_count.imm_val_reg\[23\] vssd1 vssd1 vccd1 vccd1
+ net988 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 total_design.core.regFile.register\[19\]\[1\] vssd1 vssd1 vccd1 vccd1 net2447
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09730__A1 _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 total_design.core.regFile.register\[25\]\[8\] vssd1 vssd1 vccd1 vccd1 net2458
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 total_design.core.regFile.register\[20\]\[25\] vssd1 vssd1 vccd1 vccd1 net2469
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10312__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08828_ _04048_ _04082_ _04042_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__o21ba_1
Xhold1164 total_design.keypad0.counter\[9\] vssd1 vssd1 vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07741__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1175 total_design.core.regFile.register\[30\]\[20\] vssd1 vssd1 vccd1 vccd1 net2491
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14288__Q net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1186 total_design.core.regFile.register\[17\]\[13\] vssd1 vssd1 vccd1 vccd1 net2502
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1197 total_design.core.regFile.register\[11\]\[20\] vssd1 vssd1 vccd1 vccd1 net2513
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08759_ _02918_ total_design.core.data_mem.data_cpu_i\[16\] _04013_ vssd1 vssd1 vccd1
+ vccd1 _04014_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_174_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11770_ net1742 net956 net301 _01863_ vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__a22o_1
XANTENNA__12093__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ net170 net2448 net357 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06847__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout905_X net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13440_ clknet_leaf_192_clk _00907_ net1033 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10652_ net182 net1956 net477 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__mux2_1
XANTENNA__06237__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13371_ clknet_leaf_143_clk _00838_ net1173 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10583_ net194 net1929 net369 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12322_ _01580_ _01581_ _01582_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__o21bai_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07272__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11379__A _05477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12253_ net994 _04561_ _06094_ _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__o22a_1
XFILLER_0_160_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11204_ net304 _05460_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__nand2_1
XANTENNA__07024__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12184_ total_design.core.math.pc_val\[4\] net526 _06034_ vssd1 vssd1 vccd1 vccd1
+ _01474_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11135_ _05380_ _05386_ _05388_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07980__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_X net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11066_ _05321_ _05322_ _05323_ _05324_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__or4_1
XANTENNA__10730__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10017_ net161 net2708 net416 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10222__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07732__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14198__Q net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12084__A2 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11968_ _05798_ _05825_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__nor2_4
XANTENNA__06936__A _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11652__D_N _05675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13707_ clknet_leaf_32_clk total_design.core.data_mem.stored_read_data\[14\] net1070
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[14\] sky130_fd_sc_hd__dfrtp_1
X_10919_ _05171_ _05177_ _05176_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__o21ai_1
X_11899_ _05774_ _05776_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13638_ clknet_leaf_55_clk total_design.core.data_mem.data_write_adr_i\[10\] net1117
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13569_ clknet_leaf_41_clk total_design.core.data_mem.data_bus_i\[5\] net1084 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07799__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07090_ _02633_ _02613_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__nand2b_1
XANTENNA__06671__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06471__B1 total_design.core.ctrl.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_124_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06390__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07015__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout207 _04740_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_2
X_09800_ net210 net2472 net439 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__mux2_1
Xfanout218 _04699_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
Xfanout229 net231 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__dlymetal6s2s_1
X_07992_ total_design.core.regFile.register\[25\]\[28\] net649 net591 total_design.core.regFile.register\[1\]\[28\]
+ _03488_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07971__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_163_Right_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06943_ _02493_ _02494_ net721 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_52_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09731_ net704 _04952_ _04953_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__o21ai_1
X_09662_ _04888_ _04885_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_2_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10132__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06874_ total_design.core.regFile.register\[12\]\[6\] net773 net771 total_design.core.regFile.register\[28\]\[6\]
+ _02430_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__a221o_1
XANTENNA__08110__B _03602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ _03907_ vssd1 vssd1 vccd1 vccd1 total_design.keypad0.next_rows\[3\] sky130_fd_sc_hd__inv_2
XANTENNA__09921__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09593_ net189 net2610 net455 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_141_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout266_A _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08544_ _03879_ _03882_ _03891_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__a21o_1
XANTENNA__12075__A2 _05830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08475_ total_design.keypad0.key_out\[9\] _03782_ _03810_ vssd1 vssd1 vccd1 vccd1
+ _03828_ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13740__Q total_design.core.data_bus_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07426_ total_design.core.regFile.register\[10\]\[17\] net616 net601 total_design.core.regFile.register\[31\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07357_ total_design.core.regFile.register\[26\]\[15\] net871 _02883_ _02884_ _02886_
+ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_18_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08780__B total_design.core.data_mem.data_cpu_i\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_60_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06308_ _01852_ _01881_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07254__A2 total_design.core.data_mem.data_cpu_i\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_07288_ total_design.core.regFile.register\[12\]\[14\] net774 net772 total_design.core.regFile.register\[28\]\[14\]
+ _02820_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ total_design.core.math.pc_val\[1\] net906 net755 total_design.core.data_cpu_o\[1\]
+ _04279_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06239_ _01811_ _01814_ _01817_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10307__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold250 total_design.lcd_display.row_1\[80\] vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07006__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold261 total_design.lcd_display.row_1\[109\] vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout590_X net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 total_design.lcd_display.row_1\[6\] vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold283 total_design.lcd_display.row_1\[89\] vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 total_design.lcd_display.row_2\[23\] vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout730 net731 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_2
XANTENNA__07962__B1 total_design.core.ctrl.imm_32\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout741 net743 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_165_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout752 net753 vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_4
X_09929_ net243 net2065 net425 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__mux2_1
Xfanout763 _01997_ vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__buf_4
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout774 _01994_ vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__buf_6
Xfanout785 _01986_ vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_8
Xfanout796 net797 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_4
XFILLER_0_137_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10042__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12940_ clknet_leaf_165_clk _00407_ net1158 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_161_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11510__A1 _05612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07714__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09831__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12871_ clknet_leaf_175_clk _00338_ net1052 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11822_ _05713_ _05714_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__nor2_1
XANTENNA__12066__A2 _05839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09467__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11753_ net1667 net958 net291 total_design.core.data_bus_o\[25\] vssd1 vssd1 vccd1
+ vccd1 _01381_ sky130_fd_sc_hd__a22o_1
X_14541_ net1313 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06475__B net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10704_ net236 net1930 net358 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__mux2_1
X_11684_ _05630_ net1793 net131 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14472_ clknet_leaf_40_clk _01539_ net1093 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13152__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13423_ clknet_leaf_160_clk _00890_ net1150 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10635_ net251 net2523 net478 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11601__S net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload109 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 clkload109/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13354_ clknet_leaf_25_clk _00821_ net1106 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07245__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10566_ net274 net1923 net371 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10785__C1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10725__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12305_ _06122_ _06127_ _06133_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14481__Q total_design.core.ctrl.instruction\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10217__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13285_ clknet_leaf_118_clk _00752_ net1171 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10497_ net269 net1997 net480 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12526__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12236_ net897 _06080_ net527 vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12167_ _01750_ net526 _06019_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_9_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12432__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07953__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11118_ _05365_ _05373_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__xnor2_2
X_12098_ total_design.lcd_display.row_1\[77\] _05816_ _05952_ _05954_ vssd1 vssd1
+ vccd1 vccd1 _05955_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_30_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ net352 _05240_ _05305_ _05045_ _05032_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__a32o_1
XFILLER_0_127_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11501__A1 _05679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07705__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06369__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12057__A2 _05838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06590_ total_design.core.regFile.register\[8\]\[1\] net740 net739 net723 vssd1 vssd1
+ vccd1 vccd1 _02161_ sky130_fd_sc_hd__and4_1
XANTENNA__06666__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06385__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08260_ net1388 net559 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[10\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_15_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07484__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07211_ net970 _02696_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__nand2_1
XANTENNA__06692__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08191_ total_design.core.data_mem.data_write_adr_reg\[17\] total_design.core.data_mem.data_write_adr_reg\[16\]
+ total_design.core.data_mem.data_write_adr_reg\[19\] total_design.core.data_mem.data_write_adr_reg\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__or4_1
XFILLER_0_85_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11511__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07142_ total_design.core.regFile.register\[27\]\[11\] net782 _02679_ _02680_ _02683_
+ vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_172_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07236__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07073_ total_design.core.regFile.register\[9\]\[10\] net850 net823 total_design.core.regFile.register\[19\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__a22o_1
XANTENNA__10127__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06995__A1 total_design.core.ctrl.instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_112_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07944__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07975_ total_design.core.regFile.register\[20\]\[28\] net816 _03471_ _03472_ vssd1
+ vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_143_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout383_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10801__D _05049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06926_ total_design.core.regFile.register\[10\]\[7\] net834 net798 total_design.core.regFile.register\[29\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__a22o_1
X_09714_ net466 _04898_ _04937_ _04163_ net330 vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_93_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09645_ _03465_ _04869_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__nand2b_1
X_06857_ total_design.core.regFile.register\[23\]\[6\] net680 net575 total_design.core.regFile.register\[24\]\[6\]
+ _02402_ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout648_A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09576_ _03275_ _04786_ _03326_ _03277_ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__a211o_1
XFILLER_0_171_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06788_ _02315_ _02340_ _02339_ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_69_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08527_ net932 _03863_ _03844_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_33_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08121__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout815_A _01969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ _03807_ _03811_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08791__A _02666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07409_ _02925_ _02927_ _02929_ _02935_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_137_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08389_ _03719_ _03745_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11421__S net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09098__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10420_ net185 net1974 net387 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__mux2_1
XANTENNA__07227__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10351_ net198 net2440 net489 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10037__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10782__A2 total_design.core.data_bus_o\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13070_ clknet_leaf_191_clk _00537_ net1032 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10282_ net209 net2783 net498 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout972_X net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12021_ total_design.lcd_display.row_1\[17\] _05826_ _05845_ total_design.lcd_display.row_2\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07935__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11731__B2 total_design.core.data_bus_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 _03673_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_2
Xfanout571 _02091_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__buf_4
Xfanout582 _02085_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_4
X_13972_ clknet_leaf_100_clk _01152_ net1229 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[54\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout593 net596 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__buf_6
XANTENNA__09152__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12923_ clknet_leaf_147_clk _00390_ net1152 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10500__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12039__A2 _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12854_ clknet_leaf_153_clk _00321_ net1138 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14476__Q total_design.core.ctrl.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11805_ net1863 _05704_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12785_ clknet_leaf_152_clk _00252_ net1145 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08112__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14524_ net1296 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_0_127_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11736_ net1785 net958 net290 total_design.core.data_bus_o\[8\] vssd1 vssd1 vccd1
+ vccd1 _01364_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07466__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14455_ clknet_leaf_68_clk net1404 net1109 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10295__X _05005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ _05655_ net1727 net129 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__mux2_1
X_13406_ clknet_leaf_167_clk _00873_ net1155 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10618_ net187 net2007 net366 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__mux2_1
XANTENNA__07218__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12211__A2 _02492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11598_ _05670_ net1745 net137 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__mux2_1
X_14386_ clknet_leaf_160_clk _01527_ net1142 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13337_ clknet_leaf_195_clk _00804_ net1009 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10549_ net200 total_design.core.regFile.register\[6\]\[22\] net375 vssd1 vssd1 vccd1
+ vccd1 _00829_ sky130_fd_sc_hd__mux2_1
XANTENNA__14192__RESET_B net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13268_ clknet_leaf_141_clk _00735_ net1183 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12219_ net994 _04473_ net897 vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__o21ai_1
X_13199_ clknet_leaf_146_clk _00666_ net1153 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07926__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09037__A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07760_ total_design.core.regFile.register\[20\]\[23\] net670 net612 total_design.core.regFile.register\[11\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__a22o_1
XANTENNA__08876__A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06711_ total_design.core.regFile.register\[13\]\[3\] net667 net563 total_design.core.regFile.register\[3\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__a22o_1
X_07691_ total_design.core.regFile.register\[3\]\[22\] net867 net835 total_design.core.regFile.register\[10\]\[22\]
+ _03200_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__a221o_1
XANTENNA__11506__S net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_200_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_200_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09430_ _02337_ _04104_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__or2_2
XFILLER_0_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06642_ _02211_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[2\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10410__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06396__A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09361_ _04193_ _04600_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06573_ total_design.core.regFile.register\[16\]\[1\] net854 _02125_ _02128_ _02129_
+ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_47_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08312_ net1498 net940 _03690_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[13\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11789__B2 _01795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09292_ _02689_ net504 net446 _02690_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__o22a_1
XANTENNA__07457__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08243_ net1407 net544 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[26\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_43_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09500__A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout131_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08174_ net891 _02993_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[17\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06562__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07125_ total_design.core.regFile.register\[24\]\[11\] net793 net767 total_design.core.regFile.register\[7\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08957__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1040_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1138_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07056_ total_design.core.regFile.register\[14\]\[10\] net624 net612 total_design.core.regFile.register\[11\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout598_A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout765_A _01997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ total_design.core.regFile.register\[9\]\[27\] net664 net621 total_design.core.regFile.register\[4\]\[27\]
+ _03441_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__a221o_1
X_06909_ total_design.core.regFile.register\[30\]\[7\] net662 net636 total_design.core.regFile.register\[2\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__a22o_1
X_07889_ total_design.core.regFile.register\[23\]\[26\] net811 _03376_ _03390_ vssd1
+ vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_108_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09628_ _03416_ _04188_ net505 _03417_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10320__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07696__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ _03273_ _03274_ _04186_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_3_7_0_clk_X clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_X net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12570_ net1434 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07448__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11521_ net1537 _05477_ net148 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06656__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11452_ net1802 _05651_ net157 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__mux2_1
X_14240_ clknet_leaf_109_clk _01420_ net1228 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06245__S net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10403_ net261 net2604 net386 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14171_ clknet_leaf_34_clk _01351_ net1066 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11383_ net304 _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07081__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ clknet_leaf_126_clk _00589_ net1193 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10334_ net259 net2116 net490 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13053_ clknet_leaf_11_clk _00520_ net1025 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10265_ net276 net2404 net497 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__mux2_1
XANTENNA__07908__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12004_ total_design.lcd_display.row_2\[72\] _05806_ _05834_ total_design.lcd_display.row_2\[104\]
+ _05865_ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__a221o_1
X_10196_ net2067 net390 vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout390 net393 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13955_ clknet_leaf_93_clk _01135_ net1262 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12906_ clknet_leaf_25_clk _00373_ net1106 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10230__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07687__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13886_ clknet_leaf_96_clk _01066_ net1254 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[96\]
+ sky130_fd_sc_hd__dfrtp_1
X_12837_ clknet_leaf_119_clk _00304_ net1171 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09833__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07439__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12768_ clknet_leaf_201_clk _00235_ net1004 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14507_ net72 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11640__A0 _05636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09320__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06647__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11719_ net25 net936 net879 net1839 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12699_ clknet_leaf_149_clk _00166_ net1148 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14438_ clknet_leaf_67_clk total_design.core.next_instr_wait net1112 vssd1 vssd1
+ vccd1 vccd1 total_design.core.disable_pc sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09061__A1 _04292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold805 total_design.core.regFile.register\[25\]\[18\] vssd1 vssd1 vccd1 vccd1 net2121
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14369_ clknet_leaf_106_clk _01510_ net1240 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold816 total_design.core.regFile.register\[2\]\[16\] vssd1 vssd1 vccd1 vccd1 net2132
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07072__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold827 total_design.core.regFile.register\[13\]\[21\] vssd1 vssd1 vccd1 vccd1 net2143
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 total_design.core.regFile.register\[22\]\[24\] vssd1 vssd1 vccd1 vccd1 net2154
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07611__A2 _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold849 total_design.core.regFile.register\[26\]\[17\] vssd1 vssd1 vccd1 vccd1 net2165
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09038__Y _04290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08930_ _04172_ _04183_ net316 vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10405__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08861_ total_design.core.instr_fetch _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__nor2_4
Xhold1505 total_design.core.regFile.register\[6\]\[29\] vssd1 vssd1 vccd1 vccd1 net2821
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07812_ total_design.core.regFile.register\[26\]\[24\] net645 net641 total_design.core.regFile.register\[19\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__a22o_1
Xhold1516 total_design.core.regFile.register\[27\]\[28\] vssd1 vssd1 vccd1 vccd1 net2832
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 total_design.core.regFile.register\[12\]\[6\] vssd1 vssd1 vccd1 vccd1 net2843
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08792_ total_design.core.data_mem.data_cpu_i\[8\] _02515_ vssd1 vssd1 vccd1 vccd1
+ _04047_ sky130_fd_sc_hd__and2b_1
Xhold1538 net72 vssd1 vssd1 vccd1 vccd1 net2854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1549 total_design.core.regFile.register\[20\]\[15\] vssd1 vssd1 vccd1 vccd1 net2865
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07743_ total_design.core.regFile.register\[2\]\[23\] net783 _03250_ net691 vssd1
+ vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_88_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07674_ _03184_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__inv_2
XANTENNA__10140__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09413_ total_design.core.math.pc_val\[15\] total_design.core.math.pc_val\[16\] _04609_
+ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__and3_1
X_06625_ total_design.core.regFile.register\[23\]\[2\] net810 net763 total_design.core.regFile.register\[6\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11760__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09344_ _04583_ _04584_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__or2_1
X_06556_ total_design.core.regFile.register\[29\]\[1\] net926 net946 net909 vssd1
+ vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_62_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11631__A0 _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06638__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09275_ total_design.core.data_cpu_o\[10\] net755 _04518_ net903 vssd1 vssd1 vccd1
+ vccd1 _04519_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06487_ net744 net738 net736 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__and3_4
XANTENNA_fanout513_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout134_X net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08226_ net1380 net542 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[9\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_16_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07850__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08157_ net893 _02118_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[0\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_151_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07108_ total_design.core.regFile.register\[23\]\[11\] net678 net596 total_design.core.regFile.register\[8\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__a22o_1
XANTENNA__09376__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07602__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08088_ total_design.core.regFile.register\[9\]\[30\] net665 net568 total_design.core.regFile.register\[12\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout882_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07039_ _02564_ _02584_ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06810__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10315__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ net167 total_design.core.regFile.register\[21\]\[30\] net412 vssd1 vssd1
+ vccd1 vccd1 _00357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11698__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08315__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13740_ clknet_leaf_73_clk total_design.core.data_mem.stored_write_data\[15\] net1209
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[15\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__10050__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ _05202_ _05200_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_138_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07669__A2 _03157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06467__C net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06877__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13671_ clknet_leaf_55_clk total_design.core.data_mem.data_read_adr_i\[11\] net1120
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10883_ _05140_ _05141_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_123_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12622_ clknet_leaf_186_clk _00089_ net1030 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11622__A0 _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06629__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12553_ net1486 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08094__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11504_ net1605 _05671_ net152 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__mux2_1
X_12484_ net982 net973 net884 _01696_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__a22o_1
XANTENNA__07841__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14223_ clknet_leaf_58_clk _01403_ net1126 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dfrtp_1
X_11435_ net1558 _05655_ net157 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10189__A0 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09286__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07054__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11366_ _05471_ _05476_ _05606_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__nand3_1
X_14154_ clknet_leaf_35_clk _01334_ net1068 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10733__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10317_ net202 net2143 net493 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__mux2_1
X_13105_ clknet_leaf_151_clk _00572_ net1145 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06801__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14085_ clknet_leaf_88_clk _01265_ net1260 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_11297_ _05514_ _05520_ _05554_ _05553_ _05548_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__a32o_1
XANTENNA__11689__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10248_ net219 net2227 net500 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__mux2_1
X_13036_ clknet_leaf_172_clk _00503_ net1159 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1130 net1133 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__clkbuf_2
Xfanout1141 net1144 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10179_ net189 net2721 net395 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__mux2_1
Xfanout1152 net1154 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06498__X _02072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12440__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1163 net1172 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__clkbuf_2
Xfanout1174 net1181 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__clkbuf_2
Xfanout1185 net1201 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__clkbuf_2
Xfanout1196 net1200 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_117_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13938_ clknet_leaf_85_clk _01118_ net1249 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_8__f_clk_X clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06377__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06868__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13869_ clknet_leaf_66_clk total_design.core.ctrl.imm_32\[8\] net1123 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06410_ net923 net948 net916 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__and3_2
XFILLER_0_146_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07390_ total_design.core.regFile.register\[0\]\[16\] net685 _02912_ _02916_ vssd1
+ vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__o22a_4
XANTENNA__06674__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12405__A2 _03512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11613__A0 _05645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06341_ total_design.core.ctrl.instruction\[4\] net973 vssd1 vssd1 vccd1 vccd1 _01917_
+ sky130_fd_sc_hd__nand2b_2
XFILLER_0_162_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08085__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09060_ _04158_ _04303_ _04311_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__a21oi_1
X_06272_ _01838_ _01845_ _01850_ _01836_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__and4b_1
XFILLER_0_127_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07293__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07832__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08011_ _03487_ _03506_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09034__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold602 total_design.core.regFile.register\[17\]\[0\] vssd1 vssd1 vccd1 vccd1 net1918
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold613 total_design.core.regFile.register\[5\]\[23\] vssd1 vssd1 vccd1 vccd1 net1929
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold624 total_design.core.regFile.register\[29\]\[16\] vssd1 vssd1 vccd1 vccd1 net1940
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 total_design.core.regFile.register\[25\]\[7\] vssd1 vssd1 vccd1 vccd1 net1951
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 total_design.core.regFile.register\[11\]\[30\] vssd1 vssd1 vccd1 vccd1 net1962
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 total_design.core.regFile.register\[30\]\[12\] vssd1 vssd1 vccd1 vccd1 net1973
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 total_design.core.regFile.register\[8\]\[28\] vssd1 vssd1 vccd1 vccd1 net1984
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ net254 total_design.core.regFile.register\[23\]\[10\] net418 vssd1 vssd1
+ vccd1 vccd1 _00273_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold679 total_design.core.regFile.register\[1\]\[30\] vssd1 vssd1 vccd1 vccd1 net1995
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10135__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09924__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08913_ net335 _03459_ _04166_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_110_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09893_ net250 net2568 net427 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout296_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1302 total_design.core.regFile.register\[21\]\[22\] vssd1 vssd1 vccd1 vccd1 net2618
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1313 total_design.core.regFile.register\[24\]\[15\] vssd1 vssd1 vccd1 vccd1 net2629
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08844_ net968 _01747_ _04097_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__or3_1
XANTENNA__07899__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1003_A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1324 total_design.core.regFile.register\[16\]\[27\] vssd1 vssd1 vccd1 vccd1 net2640
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1335 total_design.core.regFile.register\[29\]\[21\] vssd1 vssd1 vccd1 vccd1 net2651
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1346 total_design.core.regFile.register\[30\]\[18\] vssd1 vssd1 vccd1 vccd1 net2662
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1357 total_design.data_in_BUS\[20\] vssd1 vssd1 vccd1 vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13743__Q total_design.core.data_bus_o\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1368 total_design.core.regFile.register\[27\]\[9\] vssd1 vssd1 vccd1 vccd1 net2684
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08775_ total_design.core.data_mem.data_cpu_i\[29\] net306 _04027_ _04028_ vssd1
+ vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1379 total_design.core.regFile.register\[24\]\[13\] vssd1 vssd1 vccd1 vccd1 net2695
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06571__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07726_ net749 _03234_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[22\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06859__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07657_ total_design.core.regFile.register\[29\]\[21\] net656 net574 total_design.core.regFile.register\[24\]\[21\]
+ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout630_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout728_A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08783__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06608_ total_design.core.regFile.register\[14\]\[1\] net627 net600 total_design.core.regFile.register\[21\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07588_ total_design.core.regFile.register\[7\]\[20\] net651 net644 total_design.core.regFile.register\[26\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06539_ _02112_ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__inv_2
X_09327_ _02692_ _02743_ _02795_ _04544_ _04567_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_153_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08076__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10812__D1 _05028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09258_ _02640_ net702 _04501_ net534 vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08209_ total_design.core.data_mem.data_read_adr_reg\[9\] total_design.core.data_mem.data_read_adr_reg\[8\]
+ total_design.core.data_mem.data_read_adr_reg\[11\] total_design.core.data_mem.data_read_adr_reg\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__or4_1
X_09189_ _04336_ _04339_ net328 vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11220_ _01859_ _01869_ _01903_ _05025_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_79_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11151_ _05358_ _05399_ _05407_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__and3b_1
XANTENNA__10045__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ net225 net2579 net404 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__mux2_1
XANTENNA__09834__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11082_ _05338_ _05339_ _05340_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08958__B _02182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ net229 net2720 net410 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__mux2_1
XANTENNA__10343__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08000__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06478__B net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12096__B1 _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11984_ net474 _05831_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__nor2_4
XFILLER_0_168_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13723_ clknet_leaf_33_clk total_design.core.data_mem.stored_read_data\[30\] net1070
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[30\] sky130_fd_sc_hd__dfrtp_1
X_10935_ _05192_ _05193_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__or2_1
XANTENNA__11604__S net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ clknet_leaf_50_clk total_design.core.data_mem.data_write_adr_i\[26\] net1097
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10866_ _05102_ _05103_ _05122_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__a21bo_2
XANTENNA__06494__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10728__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14484__Q total_design.core.ctrl.instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12605_ clknet_leaf_14_clk _00072_ net1026 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08067__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13585_ clknet_leaf_37_clk total_design.core.data_mem.data_bus_i\[21\] net1076 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[21\] sky130_fd_sc_hd__dfrtp_1
X_10797_ net350 _05055_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__nor2_2
XFILLER_0_54_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07275__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12536_ net976 total_design.core.ctrl.instruction\[31\] net882 _01722_ vssd1 vssd1
+ vccd1 vccd1 _01570_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07814__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12467_ _01687_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__inv_2
XANTENNA__12435__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14206_ clknet_leaf_79_clk _01386_ net1218 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07027__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11418_ net1540 _05477_ net158 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12398_ total_design.core.math.pc_val\[28\] net989 vssd1 vssd1 vccd1 vccd1 _01657_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14137_ clknet_leaf_96_clk _01317_ net1253 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11349_ _05600_ _05602_ _05607_ _05589_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__a31o_4
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14068_ clknet_leaf_100_clk _01248_ net1229 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[86\]
+ sky130_fd_sc_hd__dfrtp_1
X_13019_ clknet_leaf_143_clk _00486_ net1173 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_06890_ total_design.core.ctrl.instruction\[25\] total_design.core.ctrl.instruction\[26\]
+ total_design.core.ctrl.instruction\[27\] vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__or3_1
XFILLER_0_146_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09045__A _04296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06388__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08560_ net1824 net338 net718 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[15\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07511_ total_design.core.regFile.register\[27\]\[18\] net779 _01992_ total_design.core.regFile.register\[20\]\[18\]
+ _03031_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__a221o_1
X_08491_ net931 total_design.keypad0.key_out\[15\] vssd1 vssd1 vccd1 vccd1 _03843_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_18_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11514__S net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07442_ total_design.core.regFile.register\[22\]\[17\] net674 net659 total_design.core.regFile.register\[30\]\[17\]
+ _02954_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07373_ total_design.core.regFile.register\[1\]\[16\] net590 net583 total_design.core.regFile.register\[6\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06324_ _01881_ _01900_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__nand2b_1
X_09112_ _04358_ _04359_ _04361_ net316 vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__o22a_1
XANTENNA__09919__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07805__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10925__Y _05184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09043_ net465 _04162_ _04294_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__o21ai_1
X_06255_ _01830_ _01833_ _01827_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__and3b_1
XFILLER_0_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11102__X _05361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07018__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold410 total_design.lcd_display.row_1\[63\] vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09558__A2 _04204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06186_ net997 _01766_ _01763_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__a21o_1
Xhold421 total_design.lcd_display.row_2\[86\] vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 net67 vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold443 total_design.lcd_display.row_2\[61\] vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold454 total_design.lcd_display.row_1\[30\] vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold465 net63 vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1120_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold476 total_design.data_in_BUS\[6\] vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold487 total_design.lcd_display.row_1\[112\] vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold498 total_design.lcd_display.row_2\[125\] vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 _02016_ vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_2
XANTENNA__07963__A _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09945_ net178 net1971 net424 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__mux2_1
Xfanout912 _01940_ vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_74_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout923 net924 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__buf_2
Xfanout934 net935 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__buf_2
Xfanout945 _03674_ vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06792__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout678_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09715__C1 _04100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout956 net959 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_146_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ net181 net2142 net431 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__mux2_1
Xfanout967 total_design.core.ctrl.instruction\[14\] vssd1 vssd1 vccd1 vccd1 net967
+ sky130_fd_sc_hd__clkbuf_4
Xfanout978 net985 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08130__Y _03622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1006_X net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1110 total_design.core.regFile.register\[24\]\[12\] vssd1 vssd1 vccd1 vccd1 net2426
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 total_design.core.program_count.imm_val_reg\[23\] vssd1 vssd1 vccd1 vccd1
+ net989 sky130_fd_sc_hd__clkbuf_2
Xhold1121 total_design.core.regFile.register\[9\]\[22\] vssd1 vssd1 vccd1 vccd1 net2437
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 total_design.core.regFile.register\[1\]\[29\] vssd1 vssd1 vccd1 vccd1 net2448
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ _04034_ _04046_ _04080_ _04081_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__and4b_1
Xhold1143 total_design.core.regFile.register\[15\]\[20\] vssd1 vssd1 vccd1 vccd1 net2459
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 total_design.core.regFile.register\[7\]\[26\] vssd1 vssd1 vccd1 vccd1 net2470
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1165 total_design.core.regFile.register\[4\]\[29\] vssd1 vssd1 vccd1 vccd1 net2481
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 total_design.core.regFile.register\[29\]\[29\] vssd1 vssd1 vccd1 vccd1 net2492
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12078__B1 _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1187 total_design.core.regFile.register\[1\]\[22\] vssd1 vssd1 vccd1 vccd1 net2503
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ _03206_ _03226_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__nand2_1
Xhold1198 total_design.core.regFile.register\[8\]\[5\] vssd1 vssd1 vccd1 vccd1 net2514
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07709_ total_design.core.regFile.register\[19\]\[22\] net641 net594 total_design.core.regFile.register\[8\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__a22o_1
X_08689_ net2522 _03957_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09494__B2 _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ net173 net2144 net360 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_172_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08049__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ net185 net2316 net477 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11372__A_N _05358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09829__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10582_ net199 total_design.core.regFile.register\[5\]\[22\] net371 vssd1 vssd1 vccd1
+ vccd1 _00861_ sky130_fd_sc_hd__mux2_1
X_13370_ clknet_leaf_132_clk _00837_ net1196 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_998 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12321_ total_design.core.math.pc_val\[20\] total_design.core.program_count.imm_val_reg\[20\]
+ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_181_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07009__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06253__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12252_ _06091_ _06093_ net994 vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12002__B1 _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06480__C net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ _05459_ _05461_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__nor2_1
X_12183_ net902 _02342_ _06033_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10564__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11134_ net515 _05048_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_196_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11065_ net520 _05044_ _05064_ _05266_ _05314_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__a32o_1
XANTENNA__10503__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ net167 net2650 net417 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14479__Q total_design.core.ctrl.instruction\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12069__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09152__X _04401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11967_ _05798_ _05809_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__nor2_4
XFILLER_0_58_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13706_ clknet_leaf_36_clk total_design.core.data_mem.stored_read_data\[13\] net1072
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[13\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10918_ _05150_ _05175_ _05168_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07496__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11898_ net35 net36 net38 net37 vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__or4b_1
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_134_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13637_ clknet_leaf_63_clk total_design.core.data_mem.data_write_adr_i\[9\] net1125
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[9\] sky130_fd_sc_hd__dfrtp_1
X_10849_ _05090_ _05093_ _05095_ _05099_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__o22ai_1
XANTENNA__07248__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13568_ clknet_leaf_41_clk total_design.core.data_mem.data_bus_i\[4\] net1092 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12519_ net975 total_design.core.instr_mem.instruction_i\[23\] vssd1 vssd1 vccd1
+ vccd1 _01714_ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06671__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13499_ clknet_leaf_149_clk _00966_ net1149 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_149_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06390__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout208 _04740_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_1
Xfanout219 _04699_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_1
X_07991_ total_design.core.regFile.register\[8\]\[28\] net594 net564 total_design.core.regFile.register\[3\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11509__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09730_ _03646_ net704 net535 vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__a21oi_1
X_06942_ total_design.core.ctrl.instruction\[28\] _02446_ vssd1 vssd1 vccd1 vccd1
+ _02494_ sky130_fd_sc_hd__nand2_1
XANTENNA__10413__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09173__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09661_ total_design.core.ctrl.instruction\[27\] net885 net755 total_design.core.data_cpu_o\[27\]
+ _04887_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__a221o_2
XFILLER_0_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06873_ total_design.core.regFile.register\[4\]\[6\] _01969_ net792 total_design.core.regFile.register\[24\]\[6\]
+ net693 vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_2_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06526__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08612_ net114 net115 net113 net112 vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__and4b_1
XANTENNA__06549__D net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09592_ _04818_ _04821_ net452 vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__a21oi_4
XANTENNA__06931__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08543_ _03879_ _03882_ _03891_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__nand3_1
XFILLER_0_65_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08474_ _03825_ _03826_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07425_ _02890_ _02940_ _02942_ _02938_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__o31a_2
XANTENNA__09228__A1 _01755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09228__B2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout426_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1168_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07239__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ total_design.core.regFile.register\[8\]\[15\] net804 _02869_ _02885_ vssd1
+ vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06307_ _01852_ _01884_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__or2_1
XANTENNA__07677__B _03187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07287_ total_design.core.regFile.register\[4\]\[14\] net815 net776 total_design.core.regFile.register\[22\]\[14\]
+ net691 vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06581__B net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06238_ net930 _01816_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__nand2_1
X_09026_ _04246_ _04278_ net449 vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout795_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06169_ total_design.core.data_cpu_o\[3\] vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__inv_2
Xhold240 total_design.lcd_display.row_1\[8\] vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 total_design.lcd_display.row_1\[31\] vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold262 total_design.lcd_display.row_1\[86\] vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold273 total_design.lcd_display.row_1\[54\] vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07411__B1 total_design.core.ctrl.imm_32\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold284 total_design.lcd_display.row_1\[11\] vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 net79 vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout962_A _01770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout583_X net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout720 _03709_ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06765__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout731 _02039_ vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_165_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09928_ net253 net2627 net422 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__mux2_1
XANTENNA__10323__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout742 net743 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__buf_1
Xfanout753 _02027_ vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__clkbuf_4
Xfanout764 _01997_ vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__clkbuf_4
Xfanout775 _01990_ vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__clkbuf_8
Xfanout786 net789 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__buf_6
Xfanout797 _01978_ vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__buf_4
X_09859_ net249 net2146 net432 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout848_X net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ clknet_leaf_197_clk _00337_ net1007 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07190__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11821_ net1878 _05711_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14540_ net1312 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XANTENNA__07478__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11752_ net1632 net958 net291 total_design.core.data_bus_o\[24\] vssd1 vssd1 vccd1
+ vccd1 _01380_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10703_ net242 net2456 net358 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__mux2_1
X_14471_ clknet_leaf_54_clk net983 net1112 vssd1 vssd1 vccd1 vccd1 total_design.core.disable_pc_reg
+ sky130_fd_sc_hd__dfrtp_1
X_11683_ _05651_ net1789 net129 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07868__A _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13422_ clknet_leaf_190_clk _00889_ net1034 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10634_ net262 net2780 net478 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13353_ clknet_leaf_177_clk _00820_ net1047 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10565_ net257 net2047 net372 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06491__B net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ _06139_ _01572_ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__nor2_1
XANTENNA__07650__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13284_ clknet_leaf_106_clk _00751_ net1233 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10496_ net276 net2439 net480 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12235_ net994 _04518_ _06078_ _06079_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11396__Y _05655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07402__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ net897 _02241_ _05758_ total_design.core.math.pc_val\[2\] _06018_ vssd1 vssd1
+ vccd1 vccd1 _06019_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_9_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10741__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06756__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11117_ _05359_ _05373_ _05374_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__or3_2
XANTENNA__10233__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ total_design.lcd_display.row_1\[45\] _05821_ _05840_ total_design.lcd_display.row_1\[53\]
+ _05953_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11048_ net352 _05210_ _05305_ _05045_ _05034_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__a32o_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07181__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09458__B2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12999_ clknet_leaf_176_clk _00466_ net1052 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06385__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07210_ net970 _02696_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08190_ total_design.core.data_mem.data_write_adr_reg\[21\] total_design.core.data_mem.data_write_adr_reg\[20\]
+ total_design.core.data_mem.data_write_adr_reg\[23\] total_design.core.data_mem.data_write_adr_reg\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__or4_1
XFILLER_0_116_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07141_ total_design.core.regFile.register\[26\]\[11\] net872 _02681_ _02682_ vssd1
+ vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10408__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07641__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07072_ total_design.core.regFile.register\[6\]\[10\] net763 net759 total_design.core.regFile.register\[21\]\[10\]
+ _02616_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_144_Left_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10528__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06747__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10143__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ total_design.core.regFile.register\[9\]\[28\] net851 net760 total_design.core.regFile.register\[21\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09932__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ net466 _04160_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__nand2_1
X_06925_ _02472_ _02474_ _02476_ _02478_ vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout376_A _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11763__A _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ _03465_ _04845_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__nor2_1
X_06856_ total_design.core.regFile.register\[6\]\[6\] net584 _02412_ net688 vssd1
+ vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07172__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_153_Left_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07305__X total_design.core.data_mem.data_cpu_i\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_96_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13751__Q total_design.core.data_bus_o\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09449__A1 _03040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09575_ net194 net2145 net453 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06787_ _02347_ vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[5\] sky130_fd_sc_hd__inv_2
XANTENNA_fanout543_A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08526_ _03861_ _03874_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08457_ _03782_ _03808_ _03810_ _03809_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout808_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08791__B net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07408_ total_design.core.regFile.register\[11\]\[16\] net795 _02931_ _02933_ _02934_
+ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_108_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07880__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08388_ _03731_ _03743_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold1560_A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07339_ total_design.core.regFile.register\[3\]\[15\] net868 net833 total_design.core.regFile.register\[31\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1240_X net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10318__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_162_Left_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10350_ net204 net2375 net489 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10782__A3 total_design.core.data_bus_o\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09009_ net472 net305 vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_167_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10281_ net216 net2415 net496 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0_clk_X clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09385__A0 _04443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ _05876_ _05877_ _05879_ _05880_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06738__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12585__RESET_B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout550 _02699_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09842__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11944__Y _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout572 _02091_ vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__buf_4
X_13971_ clknet_leaf_93_clk _01151_ net1255 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[53\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout583 _02085_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_8
Xfanout594 net596 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_171_Left_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08966__B _02868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11495__A1 _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ clknet_leaf_135_clk _00389_ net1189 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07699__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07163__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ clknet_leaf_166_clk _00320_ net1157 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06486__B net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06910__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11804_ _01729_ _05703_ _05704_ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__a21boi_1
X_12784_ clknet_leaf_186_clk _00251_ net1030 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08982__A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14523_ net1295 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
X_11735_ net1682 net958 net290 total_design.core.data_bus_o\[7\] vssd1 vssd1 vccd1
+ vccd1 _01363_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11612__S net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13373__RESET_B net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14454_ clknet_leaf_69_clk net1807 net1111 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11666_ _05679_ net1773 net130 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10736__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13405_ clknet_leaf_11_clk _00872_ net1025 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14492__Q total_design.core.ctrl.instruction\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10617_ net190 net2449 net366 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__mux2_1
XANTENNA__08415__A2 _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09612__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14385_ clknet_leaf_143_clk _01526_ net1176 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11597_ _05667_ net1641 net137 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__mux2_1
X_13336_ clknet_leaf_135_clk _00803_ net1187 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10548_ net201 net2666 net375 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_5__f_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__06977__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13267_ clknet_leaf_179_clk _00734_ net1035 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12443__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10479_ net219 net2281 net377 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__mux2_1
X_12218_ _06062_ _06063_ _06064_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13198_ clknet_leaf_189_clk _00665_ net1029 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09950__A_N total_design.core.ctrl.instruction\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__06729__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07387__C1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12149_ total_design.lcd_display.row_2\[63\] net348 _05848_ total_design.lcd_display.row_2\[127\]
+ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09128__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09752__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08876__B _02868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ total_design.core.regFile.register\[10\]\[3\] net618 net578 total_design.core.regFile.register\[27\]\[3\]
+ _02274_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__a221o_1
XANTENNA__11486__A1 _05630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07690_ total_design.core.regFile.register\[19\]\[22\] net824 net811 total_design.core.regFile.register\[23\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08595__C net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06641_ total_design.core.regFile.register\[0\]\[2\] net873 _02197_ _02210_ vssd1
+ vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_78_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06396__B _01950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06901__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09360_ _04419_ _04599_ net320 vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06572_ total_design.core.regFile.register\[22\]\[1\] net775 _02120_ _02126_ _02135_
+ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06964__X _02515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08311_ total_design.core.data_mem.data_write_adr_reg\[13\] net548 net540 total_design.core.data_mem.data_read_adr_reg\[13\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09340__X _04581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09291_ net315 _04323_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__or2_2
XFILLER_0_74_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08242_ net1439 net542 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[25\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_145_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07862__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08173_ net891 _02944_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[16\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10138__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09603__A1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07614__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07124_ total_design.core.regFile.register\[0\]\[11\] net683 _02662_ _02665_ vssd1
+ vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__o22a_4
XANTENNA__06562__D net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09927__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06968__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07055_ total_design.core.regFile.register\[23\]\[10\] net678 net616 total_design.core.regFile.register\[10\]\[10\]
+ _02599_ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1033_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14249__RESET_B net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout493_A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13746__Q total_design.core.data_bus_o\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1200_A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__A2 _01994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ total_design.core.regFile.register\[21\]\[27\] net598 _03455_ net687 vssd1
+ vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout281_X net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11477__A1 _05612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ _02455_ _02457_ _02459_ _02461_ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__or4_1
XANTENNA__10601__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ total_design.core.regFile.register\[14\]\[26\] net862 net765 total_design.core.regFile.register\[6\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__a22o_1
X_09627_ net323 _04854_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__nor2_1
X_06839_ _02028_ _02396_ total_design.core.ctrl.instruction\[26\] vssd1 vssd1 vccd1
+ vccd1 _02397_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_108_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09558_ _03282_ _04204_ _04788_ net535 vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09250__X _04495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08509_ net717 _03860_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[8\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09489_ _03137_ _04722_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11432__S net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11520_ _05674_ _05478_ _05479_ _05675_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__and4b_1
XFILLER_0_65_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07853__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07211__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11451_ net1627 _05650_ net160 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10048__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09837__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10402_ net265 net2790 net385 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__mux2_1
X_14170_ clknet_leaf_34_clk _01350_ net1066 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07605__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11382_ _05577_ _05600_ _05602_ _05607_ _05588_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__a41o_1
XFILLER_0_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06959__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13121_ clknet_leaf_123_clk _00588_ net1167 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10333_ net280 net2471 net488 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13052_ clknet_leaf_31_clk _00519_ net1061 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10264_ net246 net1837 net497 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__mux2_1
X_12003_ total_design.lcd_display.row_2\[88\] _05837_ _05848_ total_design.lcd_display.row_2\[120\]
+ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__a22o_1
XANTENNA__08030__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10195_ _04425_ net392 _04994_ vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07384__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_13__f_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout380 _05010_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11607__S net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_4
XANTENNA__11468__A1 _05679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13954_ clknet_leaf_85_clk _01134_ net1249 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10511__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07136__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ clknet_leaf_3_clk _00372_ net1012 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14487__Q total_design.core.ctrl.instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13885_ clknet_leaf_44_clk _01065_ net1089 vssd1 vssd1 vccd1 vccd1 total_design.core.mem_ctrl.next_next_data_read
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_194_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_194_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11553__D _05675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12011__B _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12836_ clknet_leaf_128_clk _00303_ net1191 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08097__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12767_ clknet_leaf_154_clk _00234_ net1136 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12438__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14506_ net72 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11718_ net23 net934 net877 net1891 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__o22a_1
XFILLER_0_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12698_ clknet_leaf_132_clk _00165_ net1196 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14437_ clknet_leaf_51_clk net1318 net1093 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_fetch
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_140_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11649_ _05650_ net1759 net135 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09597__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14368_ clknet_leaf_7_clk _01509_ net1018 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold806 total_design.core.regFile.register\[23\]\[22\] vssd1 vssd1 vccd1 vccd1 net2122
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold817 total_design.core.regFile.register\[19\]\[27\] vssd1 vssd1 vccd1 vccd1 net2133
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold828 total_design.core.regFile.register\[1\]\[28\] vssd1 vssd1 vccd1 vccd1 net2144
+ sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ clknet_leaf_172_clk _00786_ net1054 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold839 total_design.core.mem_ctrl.next_next_data_read vssd1 vssd1 vccd1 vccd1 net2155
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14299_ clknet_leaf_103_clk _00013_ net1238 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08021__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08860_ total_design.core.ctrl.instruction\[11\] net556 vssd1 vssd1 vccd1 vccd1 _04114_
+ sky130_fd_sc_hd__nand2_1
X_07811_ total_design.core.regFile.register\[16\]\[24\] net634 net602 total_design.core.regFile.register\[31\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__a22o_1
Xhold1506 total_design.core.regFile.register\[0\]\[17\] vssd1 vssd1 vccd1 vccd1 net2822
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1517 total_design.core.regFile.register\[9\]\[3\] vssd1 vssd1 vccd1 vccd1 net2833
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08791_ _02666_ net300 vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__or2_1
Xhold1528 total_design.core.regFile.register\[31\]\[14\] vssd1 vssd1 vccd1 vccd1 net2844
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 total_design.core.regFile.register\[15\]\[11\] vssd1 vssd1 vccd1 vccd1 net2855
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11517__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10421__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07742_ total_design.core.regFile.register\[5\]\[23\] net806 net759 total_design.core.regFile.register\[21\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07127__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12120__A2 _05819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07673_ _03181_ _03183_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__nor2_2
Xclkbuf_leaf_185_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_185_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09412_ _04641_ _04649_ net449 vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__a21o_1
X_06624_ total_design.core.regFile.register\[11\]\[2\] net794 net767 total_design.core.regFile.register\[7\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__a22o_1
XANTENNA__06557__D net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11760__B _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ total_design.core.math.pc_val\[12\] _04539_ total_design.core.math.pc_val\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08088__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06555_ total_design.core.regFile.register\[5\]\[1\] net921 net909 net907 vssd1 vssd1
+ vccd1 vccd1 _02128_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_158_Right_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout339_A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09274_ _04516_ _04517_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__or2_1
XANTENNA__07835__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06486_ net742 net737 net730 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08225_ net1400 net543 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[8\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_133_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1150_A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1248_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09588__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ net750 _03646_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[31\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07107_ total_design.core.regFile.register\[25\]\[11\] net650 net573 total_design.core.regFile.register\[24\]\[11\]
+ _02648_ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__a221o_1
XFILLER_0_160_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08087_ total_design.core.regFile.register\[15\]\[30\] net606 net584 total_design.core.regFile.register\[6\]\[30\]
+ _03577_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1036_X net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07038_ _02564_ _02584_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout875_A _01934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06574__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ _04240_ _04241_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__nor2_1
XANTENNA__11427__S net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10331__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12111__A2 _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10951_ _05206_ _05209_ _05057_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout830_X net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_176_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_176_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout928_X net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13670_ clknet_leaf_58_clk total_design.core.data_mem.data_read_adr_i\[10\] net1120
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[10\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06467__D net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10882_ _05118_ _05121_ _05125_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_123_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12621_ clknet_leaf_6_clk _00088_ net1017 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09421__A _02918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08079__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12552_ net1444 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06256__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08037__A _03532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06483__C net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ net1670 _05680_ net151 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12483_ net982 total_design.core.instr_mem.instruction_i\[5\] vssd1 vssd1 vccd1 vccd1
+ _01696_ sky130_fd_sc_hd__and2b_1
X_14222_ clknet_leaf_59_clk _01402_ net1126 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11434_ net1577 _05679_ net159 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__mux2_1
X_14153_ clknet_leaf_35_clk _01333_ net1068 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11365_ _05471_ _05623_ _05423_ net302 vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__o2bb2a_2
Xclkbuf_leaf_100_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10506__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13104_ clknet_leaf_182_clk _00571_ net1038 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10316_ net205 net2109 net492 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__mux2_1
X_14084_ clknet_leaf_99_clk _01264_ net1232 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11296_ _05514_ _05520_ _05554_ _05553_ _05548_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__a32oi_1
XANTENNA__11685__X _05688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08003__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13035_ clknet_leaf_114_clk _00502_ net1202 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10247_ net213 total_design.core.regFile.register\[15\]\[17\] net500 vssd1 vssd1
+ vccd1 vccd1 _00536_ sky130_fd_sc_hd__mux2_1
Xfanout1120 net1121 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__buf_2
XANTENNA__07357__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1131 net1133 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__clkbuf_4
Xfanout1142 net1144 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__clkbuf_4
X_10178_ net195 net2113 net394 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__mux2_1
Xfanout1153 net1154 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__buf_2
Xfanout1164 net1165 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__clkbuf_4
Xfanout1175 net1176 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__clkbuf_4
Xfanout1186 net1188 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10241__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08857__D net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1197 net1199 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07109__A2 _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12102__A2 _05834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13937_ clknet_leaf_94_clk _01117_ net1256 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_167_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_167_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13868_ clknet_leaf_65_clk total_design.core.ctrl.imm_32\[7\] net1123 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12819_ clknet_leaf_179_clk _00286_ net1041 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13799_ clknet_leaf_75_clk total_design.core.data_mem.data_cpu_i\[8\] net1215 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[8\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06674__B _02241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07817__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06340_ total_design.core.ctrl.instruction\[4\] net973 vssd1 vssd1 vccd1 vccd1 _01916_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09282__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10196__B net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06271_ net929 _01847_ _01849_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__and3_1
XFILLER_0_142_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08010_ _03487_ _03506_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__and2_1
XANTENNA__12617__RESET_B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold603 total_design.core.regFile.register\[4\]\[30\] vssd1 vssd1 vccd1 vccd1 net1919
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10416__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold614 total_design.core.regFile.register\[1\]\[12\] vssd1 vssd1 vccd1 vccd1 net1930
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 total_design.core.regFile.register\[27\]\[19\] vssd1 vssd1 vccd1 vccd1 net1941
+ sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap333 _02233_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold636 total_design.core.regFile.register\[24\]\[22\] vssd1 vssd1 vccd1 vccd1 net1952
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11101__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09990__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07596__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold647 total_design.core.regFile.register\[2\]\[13\] vssd1 vssd1 vccd1 vccd1 net1963
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 total_design.core.regFile.register\[10\]\[25\] vssd1 vssd1 vccd1 vccd1 net1974
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09961_ net251 net2213 net420 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__mux2_1
Xhold669 total_design.core.regFile.register\[7\]\[20\] vssd1 vssd1 vccd1 vccd1 net1985
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08912_ net471 _03415_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09892_ net261 net2458 net428 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07348__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ total_design.core.ctrl.instruction\[12\] _01746_ net967 _02029_ vssd1 vssd1
+ vccd1 vccd1 _04098_ sky130_fd_sc_hd__and4_1
Xhold1303 total_design.core.regFile.register\[12\]\[7\] vssd1 vssd1 vccd1 vccd1 net2619
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1314 total_design.core.regFile.register\[4\]\[8\] vssd1 vssd1 vccd1 vccd1 net2630
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1325 total_design.core.regFile.register\[15\]\[3\] vssd1 vssd1 vccd1 vccd1 net2641
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1336 total_design.core.regFile.register\[15\]\[12\] vssd1 vssd1 vccd1 vccd1 net2652
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10151__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1347 total_design.core.regFile.register\[31\]\[18\] vssd1 vssd1 vccd1 vccd1 net2663
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08774_ total_design.core.data_mem.data_cpu_i\[29\] net306 vssd1 vssd1 vccd1 vccd1
+ _04029_ sky130_fd_sc_hd__and2_1
Xhold1358 total_design.core.regFile.register\[23\]\[1\] vssd1 vssd1 vccd1 vccd1 net2674
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1369 total_design.core.regFile.register\[19\]\[10\] vssd1 vssd1 vccd1 vccd1 net2685
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09940__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07725_ _03229_ _03233_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_158_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_158_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout456_A _04117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07656_ total_design.core.regFile.register\[28\]\[21\] net586 net563 total_design.core.regFile.register\[3\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09241__A _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06607_ _02174_ _02175_ _02176_ _02177_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07587_ total_design.core.regFile.register\[5\]\[20\] net628 net601 total_design.core.regFile.register\[31\]\[20\]
+ _03097_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_101_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10818__C _05028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09326_ _02794_ _04565_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__nor2_1
XANTENNA__07808__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06538_ _02106_ net470 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_153_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09257_ _04499_ _04500_ net706 vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06469_ total_design.core.regFile.register\[20\]\[0\] net747 net739 net735 vssd1
+ vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08208_ total_design.core.data_mem.data_read_adr_reg\[1\] total_design.core.data_mem.data_read_adr_reg\[0\]
+ total_design.core.data_mem.data_read_adr_reg\[3\] total_design.core.data_mem.data_read_adr_reg\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09188_ _04325_ _04335_ net331 vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout992_A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11151__A_N _05358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08139_ total_design.core.regFile.register\[25\]\[31\] net648 net613 total_design.core.regFile.register\[11\]\[31\]
+ _03629_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__a221o_1
XANTENNA__10326__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07587__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ _05399_ _05407_ _05358_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__a21boi_1
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout878_X net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06795__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ net233 net2730 net405 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__mux2_1
X_11081_ net350 _05253_ _05285_ _05329_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07339__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ net238 net2331 net412 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__mux2_1
XANTENNA__09416__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10061__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09850__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__Y _05814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06478__C net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09703__X _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ net531 _05833_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__nor2_4
Xclkbuf_leaf_149_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_149_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13722_ clknet_leaf_37_clk total_design.core.data_mem.stored_read_data\[29\] net1072
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[29\] sky130_fd_sc_hd__dfrtp_1
X_10934_ _05160_ _05165_ _05167_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07511__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09151__A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13653_ clknet_leaf_51_clk total_design.core.data_mem.data_write_adr_i\[25\] net1092
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[25\] sky130_fd_sc_hd__dfrtp_1
X_10865_ _05087_ _05123_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_85_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06494__B net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12604_ clknet_leaf_30_clk _00071_ net1064 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13584_ clknet_leaf_27_clk total_design.core.data_mem.data_bus_i\[20\] net1073 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[20\] sky130_fd_sc_hd__dfrtp_1
X_10796_ _01885_ _05047_ _05053_ _05054_ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__and4_1
XFILLER_0_53_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12781__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12535_ net977 total_design.core.instr_mem.instruction_i\[31\] vssd1 vssd1 vccd1
+ vccd1 _01722_ sky130_fd_sc_hd__and2b_1
XFILLER_0_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11620__S net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12466_ total_design.keypad0.key_counter\[1\] _01686_ vssd1 vssd1 vccd1 vccd1 _01687_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10744__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14205_ clknet_leaf_110_clk _01385_ net1225 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_2
X_11417_ _05674_ _05480_ _05478_ _01855_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__and4b_2
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10236__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12397_ total_design.core.math.pc_val\[28\] net988 vssd1 vssd1 vccd1 vccd1 _01656_
+ sky130_fd_sc_hd__nand2_1
X_14136_ clknet_leaf_110_clk _01316_ net1225 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11348_ net302 _05473_ _05474_ _05606_ _05471_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__a311oi_4
X_14067_ clknet_leaf_90_clk _01247_ net1263 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12451__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ _05530_ _05537_ _05463_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__a21o_1
X_13018_ clknet_leaf_124_clk _00485_ net1188 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09724__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09760__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09613__X _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07750__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07510_ total_design.core.regFile.register\[30\]\[18\] net838 net794 total_design.core.regFile.register\[11\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08490_ net717 _03842_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[7\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_18_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07502__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07441_ total_design.core.regFile.register\[21\]\[17\] net597 net566 total_design.core.regFile.register\[12\]\[17\]
+ _02952_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06710__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07372_ total_design.core.regFile.register\[26\]\[16\] net646 net613 total_design.core.regFile.register\[11\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__a22o_1
XANTENNA__11598__A0 _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09111_ net322 _04135_ _04360_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__o21ai_1
X_06323_ _01871_ _01883_ _01900_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__or3b_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07266__A1 total_design.core.ctrl.instruction\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_128_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09042_ net466 _04167_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__nand2_1
X_06254_ net929 _01832_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08789__A_N _02868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold400 total_design.lcd_display.row_1\[120\] vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10146__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06185_ total_design.core.mem_ctrl.state\[1\] _01725_ total_design.core.mem_ctrl.state\[2\]
+ _01765_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__and4_2
XFILLER_0_130_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold411 total_design.lcd_display.row_2\[14\] vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold422 total_design.lcd_display.row_2\[93\] vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08766__A1 _03350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 total_design.lcd_display.row_2\[41\] vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09935__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold444 total_design.lcd_display.row_2\[109\] vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold455 total_design.lcd_display.row_1\[58\] vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold466 total_design.lcd_display.row_2\[28\] vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11770__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold477 total_design.lcd_display.row_2\[31\] vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11766__A _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout902 _02016_ vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__clkbuf_4
Xhold488 total_design.lcd_display.row_2\[8\] vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ net181 net2594 net423 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__mux2_1
Xhold499 total_design.lcd_display.row_2\[124\] vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 net914 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_74_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout924 _01926_ vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_4
Xfanout935 _05689_ vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__buf_2
Xfanout946 net947 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__buf_2
Xfanout957 net959 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_2
X_09875_ net187 net2278 net431 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__mux2_1
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout968 net970 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__clkbuf_4
Xhold1100 total_design.core.regFile.register\[14\]\[31\] vssd1 vssd1 vccd1 vccd1 net2416
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13754__Q total_design.core.data_bus_o\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout573_A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout979 net985 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__buf_2
Xhold1111 total_design.core.regFile.register\[8\]\[30\] vssd1 vssd1 vccd1 vccd1 net2427
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1122 total_design.core.regFile.register\[8\]\[21\] vssd1 vssd1 vccd1 vccd1 net2438
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ _02613_ net310 _04043_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__or3_1
Xhold1133 total_design.core.regFile.register\[4\]\[24\] vssd1 vssd1 vccd1 vccd1 net2449
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 total_design.core.regFile.register\[8\]\[25\] vssd1 vssd1 vccd1 vccd1 net2460
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 total_design.core.regFile.register\[12\]\[4\] vssd1 vssd1 vccd1 vccd1 net2471
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07741__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1166 total_design.core.regFile.register\[25\]\[1\] vssd1 vssd1 vccd1 vccd1 net2482
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1177 total_design.core.regFile.register\[13\]\[11\] vssd1 vssd1 vccd1 vccd1 net2493
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ _03253_ _03273_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__and2_1
Xhold1188 total_design.core.regFile.register\[22\]\[23\] vssd1 vssd1 vccd1 vccd1 net2504
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout740_A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1199 total_design.core.regFile.register\[21\]\[28\] vssd1 vssd1 vccd1 vccd1 net2515
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__B _02818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07708_ total_design.core.regFile.register\[26\]\[22\] net645 net590 total_design.core.regFile.register\[1\]\[22\]
+ _03216_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__a221o_1
X_08688_ _03959_ _03962_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ total_design.core.regFile.register\[3\]\[21\] net867 net760 total_design.core.regFile.register\[21\]\[21\]
+ _03150_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10650_ net189 net2766 net477 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11589__A0 _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09309_ _04460_ _04550_ net326 vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__mux2_1
X_10581_ net201 net2451 net371 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11440__S net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12320_ total_design.core.math.pc_val\[19\] net522 _01586_ _01587_ vssd1 vssd1 vccd1
+ vccd1 _01489_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11012__Y _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12251_ _06082_ _06083_ _06084_ _06092_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_146_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10056__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09403__C1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11379__C _05626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11202_ _05460_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__inv_2
XANTENNA__09845__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12182_ net898 _06031_ _06032_ net526 vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__a31o_1
XANTENNA__06768__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08969__B _02818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ net511 _05047_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__nor2_2
XANTENNA__07873__B _03375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07980__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ _05045_ _05078_ _05268_ _05314_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__a22o_1
XANTENNA__06489__B net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ net171 net2167 net414 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__mux2_1
XANTENNA__07193__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07732__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output123_A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11615__S net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11966_ total_design.lcd_display.row_1\[16\] _05826_ _05827_ total_design.lcd_display.row_1\[32\]
+ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__a22o_1
XANTENNA__10739__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10917_ _05150_ _05168_ _05171_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__or3b_1
XFILLER_0_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ clknet_leaf_37_clk total_design.core.data_mem.stored_read_data\[12\] net1076
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11897_ net35 net36 net38 net37 vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13636_ clknet_leaf_66_clk total_design.core.data_mem.data_write_adr_i\[8\] net1122
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[8\] sky130_fd_sc_hd__dfrtp_1
X_10848_ _05105_ _05106_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09237__A2 _02565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13567_ clknet_leaf_41_clk total_design.core.data_mem.data_bus_i\[3\] net1090 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12446__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10779_ total_design.core.data_bus_o\[19\] total_design.core.data_bus_o\[22\] total_design.core.data_bus_o\[28\]
+ total_design.core.data_bus_o\[30\] net696 vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__o41a_1
XFILLER_0_55_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07799__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12518_ net976 net966 net881 _01713_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13498_ clknet_leaf_124_clk _00965_ net1187 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12449_ net2663 net216 net344 vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09755__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__B2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06759__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08879__B _02770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11586__A _05478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14119_ clknet_leaf_84_clk _01299_ net1243 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_35_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07990_ net554 _03486_ _03179_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__a21oi_1
Xfanout209 _04721_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_157_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07971__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06941_ total_design.core.ctrl.instruction\[28\] _02446_ vssd1 vssd1 vccd1 vccd1
+ _02493_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_52_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09660_ net904 _04886_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06872_ total_design.core.regFile.register\[5\]\[6\] net807 _02425_ _02427_ _02428_
+ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_2_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07184__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08611_ net112 net114 net115 net113 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.next_rows\[1\]
+ sky130_fd_sc_hd__nand4b_2
XFILLER_0_94_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09591_ net903 _04819_ _04820_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11525__S net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08542_ _03889_ _03890_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08473_ _03798_ _03824_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout154_A _05681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07424_ _02948_ vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[17\] sky130_fd_sc_hd__inv_2
XANTENNA__09228__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07355_ total_design.core.regFile.register\[17\]\[15\] net821 net817 total_design.core.regFile.register\[20\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout419_A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06306_ _01852_ _01884_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07286_ total_design.core.regFile.register\[26\]\[14\] net869 net779 total_design.core.regFile.register\[27\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13749__Q total_design.core.data_bus_o\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06998__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09025_ _02338_ _04277_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__nand2_1
X_06237_ total_design.core.data_adr_o\[21\] _01815_ net961 vssd1 vssd1 vccd1 vccd1
+ _01816_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1230_A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold230 total_design.lcd_display.row_1\[46\] vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 total_design.lcd_display.row_1\[21\] vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
X_06168_ total_design.core.math.pc_val\[2\] vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_148_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold252 total_design.lcd_display.row_1\[32\] vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 total_design.lcd_display.row_1\[56\] vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08789__B total_design.core.data_mem.data_cpu_i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold274 total_design.lcd_display.row_1\[18\] vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07411__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold285 net125 vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10604__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold296 total_design.lcd_display.row_1\[35\] vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 _03927_ vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__buf_2
Xfanout721 _02150_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__buf_2
XANTENNA__07962__A2 total_design.core.data_mem.data_cpu_i\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout732 net733 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09927_ net250 net2013 net424 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout743 _02031_ vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_2
XANTENNA_fanout955_A _01911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout576_X net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout754 net755 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_4
Xfanout765 _01997_ vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_8
Xfanout776 _01990_ vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_2
Xfanout787 net789 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_8
X_09858_ net261 net2221 net432 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout798 net801 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__buf_6
XANTENNA__07714__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08809_ net311 total_design.core.data_mem.data_cpu_i\[6\] vssd1 vssd1 vccd1 vccd1
+ _04064_ sky130_fd_sc_hd__nand2_1
X_09789_ net263 net2804 net440 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13861__D total_design.core.ctrl.imm_32\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06922__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11435__S net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11820_ total_design.lcd_display.cnt_20ms\[12\] _05711_ vssd1 vssd1 vccd1 vccd1 _05713_
+ sky130_fd_sc_hd__and2_1
X_11751_ net1648 net958 net292 total_design.core.data_bus_o\[23\] vssd1 vssd1 vccd1
+ vccd1 _01379_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout910_X net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_80_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10702_ net255 net2285 net357 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__mux2_1
X_14470_ clknet_leaf_54_clk net1383 net1110 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11682_ _05650_ net1697 net130 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13421_ clknet_leaf_1_clk _00888_ net1005 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10633_ _04452_ net1944 net476 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10234__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13352_ clknet_leaf_171_clk _00819_ net1056 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10564_ net281 net2856 net369 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__mux2_1
XANTENNA__10785__A1 total_design.core.data_bus_o\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ total_design.core.math.pc_val\[18\] total_design.core.program_count.imm_val_reg\[18\]
+ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06491__C net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13283_ clknet_leaf_5_clk _00750_ net1023 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10495_ net246 net1897 net481 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09575__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12234_ _06076_ _06077_ net994 vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12526__A2 total_design.core.ctrl.instruction\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12165_ _05760_ _06014_ _06015_ net526 vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__a31oi_1
XANTENNA__10514__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ _05373_ _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__nor2_1
XANTENNA__07953__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12096_ total_design.lcd_display.row_1\[5\] _05830_ _05849_ total_design.lcd_display.row_2\[53\]
+ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__a22o_1
XANTENNA__09155__A1 _02367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11047_ net352 _05208_ _05305_ _05045_ _05031_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_30_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07166__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07705__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
X_12998_ clknet_leaf_200_clk _00465_ net1001 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11949_ _05732_ _05742_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__nand2b_4
Xclkbuf_leaf_71_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08130__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10473__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13619_ clknet_leaf_49_clk net1323 net1102 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06692__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07140_ total_design.core.regFile.register\[16\]\[11\] net854 net797 total_design.core.regFile.register\[11\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07071_ total_design.core.regFile.register\[25\]\[10\] net842 net806 total_design.core.regFile.register\[5\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10424__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07944__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07973_ total_design.core.regFile.register\[16\]\[28\] net855 net811 total_design.core.regFile.register\[23\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_143_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09712_ net332 _04854_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__or2_1
X_06924_ total_design.core.regFile.register\[13\]\[7\] net789 net758 total_design.core.regFile.register\[4\]\[7\]
+ _02477_ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__a221o_1
XANTENNA__09146__B2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12150__B1 _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ _04869_ _03465_ _04845_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__and3b_1
X_06855_ total_design.core.regFile.register\[5\]\[6\] net630 net626 total_design.core.regFile.register\[14\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout271_A _04348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06904__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout369_A _05013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09574_ net506 _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__and2_1
X_06786_ net721 _02345_ _02346_ _02344_ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__o211a_2
XANTENNA_clkbuf_leaf_180_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08525_ _03864_ _03874_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_69_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1180_A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout157_X net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08121__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ total_design.keypad0.key_out\[8\] net933 vssd1 vssd1 vccd1 vccd1 _03810_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_0_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07407_ total_design.core.regFile.register\[9\]\[16\] net852 net800 total_design.core.regFile.register\[29\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08387_ _03731_ _03743_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__and2_1
XANTENNA__06683__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_195_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout703_A _04204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10216__A0 _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07338_ _02853_ _02854_ _02867_ net685 total_design.core.regFile.register\[0\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__o32a_4
XFILLER_0_144_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13672__RESET_B net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07269_ total_design.core.regFile.register\[9\]\[14\] _02049_ net633 total_design.core.regFile.register\[16\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_115_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12508__A2 total_design.core.ctrl.instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09008_ net331 _04252_ _04260_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_167_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10782__A4 total_design.core.data_bus_o\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10280_ net215 net2039 net496 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10334__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12115__A _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07396__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07935__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07209__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_133_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 _03676_ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09137__A1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout551 _02108_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__buf_4
Xfanout562 net565 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_8
X_13970_ clknet_leaf_86_clk _01150_ net1247 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[52\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout573 net576 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_8
Xfanout584 _02085_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12141__B1 _05840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_4
X_12921_ clknet_leaf_188_clk _00388_ net1029 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09143__B _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_148_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12852_ clknet_leaf_142_clk _00319_ net1182 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06486__C net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11803_ total_design.lcd_display.cnt_20ms\[4\] _03911_ vssd1 vssd1 vccd1 vccd1 _05704_
+ sky130_fd_sc_hd__nand2_1
X_12783_ clknet_leaf_146_clk _00250_ net1178 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08982__B _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08112__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14522_ net1294 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
X_11734_ net1810 net957 net290 total_design.core.data_bus_o\[6\] vssd1 vssd1 vccd1
+ vccd1 _01362_ sky130_fd_sc_hd__a22o_1
XANTENNA__06783__A total_design.core.ctrl.instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07320__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11665_ _05632_ net1734 net131 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__mux2_1
X_14453_ clknet_leaf_67_clk net1373 net1111 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10509__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10207__A0 _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10616_ net193 net2368 net365 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__mux2_1
X_13404_ clknet_leaf_28_clk _00871_ net1075 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14384_ clknet_leaf_179_clk _01525_ net1041 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11596_ _05665_ net1769 net138 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07084__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13335_ clknet_leaf_161_clk _00802_ net1151 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06426__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10547_ net207 net2140 net373 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13266_ clknet_leaf_138_clk _00733_ net1185 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10478_ net214 net2355 net377 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10752__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12217_ _06062_ _06063_ net995 vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10244__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13197_ clknet_leaf_7_clk _00664_ net1016 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07926__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ total_design.lcd_display.row_1\[111\] _05829_ _05971_ _06002_ vssd1 vssd1
+ vccd1 vccd1 _06003_ sky130_fd_sc_hd__a211o_1
X_12079_ total_design.lcd_display.row_1\[124\] _05843_ _05846_ total_design.lcd_display.row_2\[100\]
+ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07139__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06640_ _02199_ _02203_ _02206_ _02209_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__or4_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12435__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06571_ total_design.core.regFile.register\[19\]\[1\] net823 net793 total_design.core.regFile.register\[24\]\[1\]
+ _02143_ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_44_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08892__B _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08310_ net1481 net940 _03689_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[12\]
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_47_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09290_ net319 _04337_ net295 vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ net1474 net543 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[24\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_157_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06665__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10419__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08172_ net892 _02893_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[15\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_136_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07123_ _02649_ _02653_ _02654_ _02664_ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__or4_1
XFILLER_0_160_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07054_ total_design.core.regFile.register\[26\]\[10\] net644 net573 total_design.core.regFile.register\[24\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__a22o_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__clkbuf_4
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07378__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1026_A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09943__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09119__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_A _05007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09119__B2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ total_design.core.regFile.register\[30\]\[27\] net660 net637 total_design.core.regFile.register\[2\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__a22o_1
XANTENNA__12123__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06907_ total_design.core.regFile.register\[7\]\[7\] net652 net632 total_design.core.regFile.register\[16\]\[7\]
+ _02460_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a221o_1
X_07887_ total_design.core.regFile.register\[26\]\[26\] net870 net807 total_design.core.regFile.register\[5\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout653_A _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06838_ _02149_ _02345_ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__and2_1
X_09626_ net465 _04852_ _04851_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_108_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07550__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09557_ net705 _04787_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__nor2_1
X_06769_ total_design.core.regFile.register\[30\]\[4\] net659 _02330_ net686 vssd1
+ vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout820_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout918_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ total_design.data_in_BUS\[8\] net342 _03859_ vssd1 vssd1 vccd1 vccd1 _03860_
+ sky130_fd_sc_hd__a21oi_1
X_09488_ _03086_ _04701_ _03085_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07302__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08439_ _03792_ _03793_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_92_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06656__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10329__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11450_ net1801 _05633_ net159 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10401_ net274 net2372 net386 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11381_ net304 net510 _05034_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__or3b_1
XFILLER_0_116_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13120_ clknet_leaf_193_clk _00587_ net1012 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10332_ net269 net2444 net488 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__mux2_1
XANTENNA__07081__A2 _01992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09419__A _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13051_ clknet_leaf_147_clk _00518_ net1152 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10064__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10263_ net286 net2835 net497 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__mux2_1
X_12002_ total_design.lcd_display.row_2\[64\] _05819_ _05853_ total_design.lcd_display.row_2\[112\]
+ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a221o_1
XANTENNA__07908__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09853__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ net2135 net393 vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout370 _05013_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout381 net384 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_6
Xfanout392 net393 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_8
X_13953_ clknet_leaf_94_clk _01133_ net1256 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_21_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12904_ clknet_leaf_24_clk _00371_ net1055 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13884_ clknet_leaf_39_clk total_design.core.ctrl.imm_32\[23\] net1095 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[23\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07541__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12835_ clknet_leaf_16_clk _00302_ net1022 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_26_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11623__S net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12766_ clknet_leaf_174_clk _00233_ net1155 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10747__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14505_ clknet_leaf_51_clk _00003_ net1092 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instr_fetch
+ sky130_fd_sc_hd__dfrtp_1
X_11717_ net22 net934 net877 net1739 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__o22a_1
XANTENNA__06647__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12697_ clknet_leaf_194_clk _00164_ net1010 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10239__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11648_ _05633_ net1696 net135 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__mux2_1
X_14436_ clknet_leaf_37_clk total_design.core.data_out_INSTR\[31\] net1076 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[31\] sky130_fd_sc_hd__dfrtp_1
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 en vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_1
X_11579_ _05643_ net1597 net141 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__mux2_1
XANTENNA__12454__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14367_ clknet_leaf_126_clk _01508_ net1193 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold807 total_design.core.regFile.register\[20\]\[6\] vssd1 vssd1 vccd1 vccd1 net2123
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13318_ clknet_leaf_197_clk _00785_ net1007 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07072__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold818 total_design.core.regFile.register\[30\]\[13\] vssd1 vssd1 vccd1 vccd1 net2134
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold829 total_design.core.regFile.register\[30\]\[23\] vssd1 vssd1 vccd1 vccd1 net2145
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ clknet_leaf_102_clk _00012_ net1238 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13249_ clknet_leaf_118_clk _00716_ net1169 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09763__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07810_ total_design.core.regFile.register\[22\]\[24\] net675 net664 total_design.core.regFile.register\[9\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__a22o_1
XANTENNA__10702__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1507 total_design.core.regFile.register\[25\]\[12\] vssd1 vssd1 vccd1 vccd1 net2823
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08790_ total_design.core.data_mem.data_cpu_i\[15\] _02868_ vssd1 vssd1 vccd1 vccd1
+ _04045_ sky130_fd_sc_hd__and2b_1
Xhold1518 total_design.core.regFile.register\[28\]\[22\] vssd1 vssd1 vccd1 vccd1 net2834
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12105__B1 _05850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08309__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1529 total_design.core.instr_mem.instruction_i\[3\] vssd1 vssd1 vccd1 vccd1 net2845
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07780__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ total_design.core.regFile.register\[16\]\[23\] net854 net838 total_design.core.regFile.register\[30\]\[23\]
+ _03237_ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_88_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08324__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07672_ net299 _03180_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09411_ _04642_ _04643_ _04648_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__and3_1
X_06623_ total_design.core.regFile.register\[18\]\[2\] net860 net779 total_design.core.regFile.register\[27\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_17_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11533__S net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ total_design.core.math.pc_val\[12\] total_design.core.math.pc_val\[13\] _04539_
+ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_138_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06554_ total_design.core.regFile.register\[8\]\[1\] net920 net919 net913 vssd1 vssd1
+ vccd1 vccd1 _02127_ sky130_fd_sc_hd__and4_1
XFILLER_0_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09273_ total_design.core.math.pc_val\[9\] _04471_ total_design.core.math.pc_val\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06638__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10149__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06485_ total_design.core.regFile.register\[19\]\[0\] net747 net737 net733 vssd1
+ vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__and4_1
XFILLER_0_114_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08224_ net1356 net545 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[7\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09938__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08155_ _03623_ _03645_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_31_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout401_A _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07599__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1143_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07106_ total_design.core.regFile.register\[20\]\[11\] net673 net582 total_design.core.regFile.register\[6\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__a22o_1
XANTENNA__07063__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08086_ total_design.core.regFile.register\[13\]\[30\] net668 net564 total_design.core.regFile.register\[3\]\[30\]
+ _03578_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07037_ net552 total_design.core.data_mem.data_cpu_i\[9\] total_design.core.ctrl.imm_32\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a21o_1
XANTENNA__06810__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09526__X _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_X net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A _01941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10612__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ net469 net311 vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07939_ _03431_ _03433_ _03438_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout656_X net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08315__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10950_ _05203_ _05205_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_127_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09609_ total_design.core.math.pc_val\[24\] total_design.core.math.pc_val\[25\] _04799_
+ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_27_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10881_ _05121_ _05125_ _05118_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__a21boi_2
XANTENNA__06877__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11443__S net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12620_ clknet_leaf_169_clk _00087_ net1159 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09276__B1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06537__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12551_ net1426 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06629__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07287__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10059__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ net1546 _05655_ net149 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12482_ net980 total_design.core.ctrl.instruction\[4\] net884 _01695_ vssd1 vssd1
+ vccd1 vccd1 _01543_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09579__A1 _03329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14221_ clknet_leaf_57_clk _01401_ net1115 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dfrtp_1
X_11433_ net302 _05653_ _05658_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_163_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14152_ clknet_leaf_35_clk _01332_ net1068 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11364_ _05476_ _05606_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__xor2_1
XANTENNA__07054__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13103_ clknet_leaf_147_clk _00570_ net1150 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10315_ net212 net2422 net493 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__mux2_1
X_14083_ clknet_leaf_89_clk _01263_ net1260 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06801__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11295_ _05515_ _05551_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__xor2_2
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13034_ clknet_leaf_25_clk _00501_ net1106 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10246_ net220 net2339 net502 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__mux2_1
XANTENNA__11689__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09200__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1110 net1121 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__buf_2
Xfanout1121 net1134 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__buf_2
XANTENNA__11618__S net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1132 net1133 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__buf_2
X_10177_ net197 net2157 net395 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__mux2_1
XANTENNA__10522__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1143 net1144 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07762__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1154 net1172 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__clkbuf_2
Xfanout1165 net1168 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14498__Q total_design.core.ctrl.instruction\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1176 net1181 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06301__A _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1187 net1188 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__clkbuf_2
Xfanout1198 net1199 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08306__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13936_ clknet_leaf_98_clk _01116_ net1241 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06868__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13867_ clknet_leaf_65_clk total_design.core.ctrl.imm_32\[6\] net1124 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12449__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12818_ clknet_leaf_145_clk _00285_ net1179 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09267__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13798_ clknet_leaf_76_clk total_design.core.data_mem.data_cpu_i\[7\] net1213 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12749_ clknet_leaf_4_clk _00216_ net1023 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09758__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06270_ total_design.core.data_adr_o\[10\] _01848_ net963 vssd1 vssd1 vccd1 vccd1
+ _01849_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07293__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14419_ clknet_leaf_32_clk total_design.core.data_out_INSTR\[14\] net1062 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[14\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11377__A1 total_design.core.data_bus_o\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold604 total_design.core.regFile.register\[22\]\[1\] vssd1 vssd1 vccd1 vccd1 net1920
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold615 total_design.core.regFile.register\[18\]\[11\] vssd1 vssd1 vccd1 vccd1 net1931
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 total_design.core.regFile.register\[18\]\[26\] vssd1 vssd1 vccd1 vccd1 net1942
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold637 total_design.core.regFile.register\[20\]\[2\] vssd1 vssd1 vccd1 vccd1 net1953
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold648 total_design.core.regFile.register\[17\]\[30\] vssd1 vssd1 vccd1 vccd1 net1964
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 total_design.core.regFile.register\[25\]\[21\] vssd1 vssd1 vccd1 vccd1 net1975
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ net261 net2723 net420 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire457_X net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08911_ _04164_ _04162_ net465 vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09891_ net267 net1951 net426 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__mux2_1
XANTENNA__11528__S net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10432__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09813__A_N total_design.core.ctrl.instruction\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08842_ total_design.core.ctrl.instruction\[12\] _02029_ vssd1 vssd1 vccd1 vccd1
+ _04097_ sky130_fd_sc_hd__nand2_1
Xhold1304 total_design.core.regFile.register\[25\]\[29\] vssd1 vssd1 vccd1 vccd1 net2620
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07753__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1315 total_design.core.regFile.register\[23\]\[29\] vssd1 vssd1 vccd1 vccd1 net2631
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1326 total_design.core.regFile.register\[24\]\[23\] vssd1 vssd1 vccd1 vccd1 net2642
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1337 total_design.core.regFile.register\[12\]\[17\] vssd1 vssd1 vccd1 vccd1 net2653
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08773_ _03486_ _03506_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__or2_1
Xhold1348 total_design.core.regFile.register\[1\]\[14\] vssd1 vssd1 vccd1 vccd1 net2664
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 total_design.core.regFile.register\[13\]\[18\] vssd1 vssd1 vccd1 vccd1 net2675
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07724_ _03183_ _03232_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__nor2_2
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07505__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07655_ total_design.core.regFile.register\[20\]\[21\] net671 net571 total_design.core.regFile.register\[17\]\[21\]
+ _03163_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__a221o_1
XANTENNA__06859__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06606_ total_design.core.regFile.register\[10\]\[1\] net616 _02154_ _02159_ _02166_
+ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout449_A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07313__Y _02845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07586_ total_design.core.regFile.register\[22\]\[20\] net674 net659 total_design.core.regFile.register\[30\]\[20\]
+ _03094_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09325_ _02743_ _04545_ _02795_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06584__C net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06537_ total_design.core.data_mem.data_cpu_i\[0\] total_design.core.ctrl.imm_32\[0\]
+ net551 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout616_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10812__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ _02637_ _04498_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_10__f_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06468_ net744 net738 net734 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08207_ total_design.core.data_mem.data_read_adr_reg\[5\] total_design.core.data_mem.data_read_adr_reg\[4\]
+ total_design.core.data_mem.data_read_adr_reg\[7\] total_design.core.data_mem.data_read_adr_reg\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09187_ _04432_ _04433_ net319 vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06399_ total_design.core.regFile.register\[8\]\[0\] net922 net919 net913 vssd1 vssd1
+ vccd1 vccd1 _01975_ sky130_fd_sc_hd__and4_1
XANTENNA__10607__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08138_ total_design.core.regFile.register\[20\]\[31\] net671 net602 total_design.core.regFile.register\[31\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07036__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08069_ total_design.core.regFile.register\[1\]\[30\] net829 net804 total_design.core.regFile.register\[8\]\[30\]
+ _03560_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__a221o_1
XANTENNA__07992__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ net228 net2333 net405 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__mux2_1
X_11080_ net350 _05280_ _05290_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11438__S net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ net242 net2655 net413 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__mux2_1
XANTENNA__10342__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11540__A1 _05652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12096__A2 _05830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11982_ net531 _05817_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__nor2_4
X_13721_ clknet_leaf_35_clk total_design.core.data_mem.stored_read_data\[28\] net1071
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10933_ _05165_ _05167_ _05160_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06267__S net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13652_ clknet_leaf_50_clk total_design.core.data_mem.data_write_adr_i\[24\] net1097
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10864_ _05122_ _05121_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12603_ clknet_leaf_150_clk _00070_ net1173 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10795_ total_design.core.data_bus_o\[14\] net698 vssd1 vssd1 vccd1 vccd1 _05054_
+ sky130_fd_sc_hd__nand2_1
X_13583_ clknet_leaf_37_clk total_design.core.data_mem.data_bus_i\[19\] net1076 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07275__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12534_ net974 total_design.core.ctrl.instruction\[30\] net881 _01721_ vssd1 vssd1
+ vccd1 vccd1 _01569_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07680__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12465_ net1887 _05785_ _01686_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10517__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14204_ clknet_leaf_80_clk _01384_ net1222 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11416_ _01859_ _01861_ _01869_ _01903_ _01854_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a2111o_2
XANTENNA__07027__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12396_ total_design.core.math.pc_val\[27\] net523 _01654_ _01655_ vssd1 vssd1 vccd1
+ vccd1 _01497_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08214__C _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11347_ _05462_ _05604_ _05605_ _05470_ _05440_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__a32o_2
X_14135_ clknet_leaf_83_clk _01315_ net1243 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07893__Y _03395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08775__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07983__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14066_ clknet_leaf_88_clk _01246_ net1250 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[84\]
+ sky130_fd_sc_hd__dfrtp_1
X_11278_ _05442_ _05447_ _05535_ _05533_ _05532_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__a32o_1
XANTENNA__09724__A1 total_design.core.ctrl.instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13017_ clknet_leaf_196_clk _00484_ net1028 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10229_ _04113_ _04972_ _05002_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__or3_1
XANTENNA__09724__B2 total_design.core.data_cpu_o\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10252__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11531__A1 _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__B net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 total_design.core.data_mem.data_cpu_i_reg\[6\] vssd1 vssd1 vccd1 vccd1 net1317
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_146_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13919_ clknet_leaf_97_clk _01099_ net1244 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07440_ total_design.core.regFile.register\[15\]\[17\] net604 _02963_ net686 vssd1
+ vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07371_ total_design.core.regFile.register\[9\]\[16\] net665 net599 total_design.core.regFile.register\[21\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09110_ net324 _04182_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__or2_1
X_06322_ _01871_ _01883_ _01900_ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07797__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09041_ net465 _04164_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__nand2_1
XANTENNA__06474__B1 total_design.core.ctrl.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_06253_ total_design.core.data_adr_o\[22\] _01831_ net961 vssd1 vssd1 vccd1 vccd1
+ _01832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07018__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06184_ _01764_ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__inv_2
Xhold401 total_design.lcd_display.row_2\[81\] vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09412__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold412 total_design.core.math.pc_val\[4\] vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 total_design.data_in_BUS\[28\] vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 net61 vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08766__A2 _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold445 total_design.lcd_display.row_1\[4\] vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold456 total_design.lcd_display.row_2\[113\] vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold467 total_design.keypad0.counter\[8\] vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07974__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold478 total_design.lcd_display.row_1\[19\] vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11766__B _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold489 total_design.lcd_display.row_2\[115\] vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09943_ net187 net1970 net423 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout903 net904 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__buf_4
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout914 net915 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout925 _01925_ vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__clkbuf_2
Xfanout936 _05688_ vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout399_A _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10162__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ net191 net2596 net431 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__mux2_1
Xfanout947 _01942_ vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__buf_2
Xfanout958 net959 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_146_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout969 net970 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__clkbuf_2
Xhold1101 total_design.core.regFile.register\[12\]\[27\] vssd1 vssd1 vccd1 vccd1 net2417
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1106_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1112 total_design.core.regFile.register\[10\]\[23\] vssd1 vssd1 vccd1 vccd1 net2428
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1123 total_design.core.regFile.register\[7\]\[2\] vssd1 vssd1 vccd1 vccd1 net2439
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ _04037_ _04041_ _04055_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__or3_1
Xhold1134 total_design.core.regFile.register\[24\]\[29\] vssd1 vssd1 vccd1 vccd1 net2450
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 total_design.core.regFile.register\[15\]\[19\] vssd1 vssd1 vccd1 vccd1 net2461
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A _02092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1156 total_design.core.regFile.register\[28\]\[19\] vssd1 vssd1 vccd1 vccd1 net2472
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 total_design.core.regFile.register\[21\]\[9\] vssd1 vssd1 vccd1 vccd1 net2483
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12078__A2 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09479__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1178 total_design.core.regFile.register\[3\]\[0\] vssd1 vssd1 vccd1 vccd1 net2494
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ _03253_ _03273_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__nor2_1
Xhold1189 total_design.core.regFile.register\[19\]\[2\] vssd1 vssd1 vccd1 vccd1 net2505
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_136_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07707_ total_design.core.regFile.register\[29\]\[22\] net656 net567 total_design.core.regFile.register\[12\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08687_ total_design.keypad0.counter\[16\] _03958_ vssd1 vssd1 vccd1 vccd1 _03962_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_67_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout354_X net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ total_design.core.regFile.register\[9\]\[21\] net852 net768 total_design.core.regFile.register\[7\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_172_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07569_ _03064_ _03084_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09398__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09308_ _04504_ _04549_ net460 vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__mux2_1
X_10580_ net206 net2611 net369 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10337__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09239_ _04390_ _04483_ net326 vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_9__f_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12250_ _06082_ _06083_ _06084_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_118_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07009__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12002__A2 _05819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11201_ net515 _05047_ _05053_ _05054_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__nand4_2
X_12181_ net994 _04371_ _04372_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ _05385_ _05388_ _05390_ _05379_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__o22ai_4
Xhold990 total_design.core.regFile.register\[27\]\[20\] vssd1 vssd1 vccd1 vccd1 net2306
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11063_ net350 net180 _05045_ _05035_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10072__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11513__A1 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ net174 net2872 net416 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__mux2_1
XANTENNA__09861__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06489__C net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08985__B _02515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12069__A2 _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07234__X _02770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11965_ _05807_ _05820_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__nor2_4
XFILLER_0_99_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08142__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ clknet_leaf_38_clk total_design.core.data_mem.stored_read_data\[11\] net1078
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[11\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ _05165_ _05167_ _05171_ _05172_ _05173_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_80_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07496__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ net35 net36 net37 net38 vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__or4b_2
XFILLER_0_86_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13635_ clknet_leaf_60_clk total_design.core.data_mem.data_write_adr_i\[7\] net1131
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[7\] sky130_fd_sc_hd__dfrtp_1
X_10847_ _05099_ _05100_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07248__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13566_ clknet_leaf_41_clk total_design.core.data_mem.data_bus_i\[2\] net1092 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10778_ net1266 total_design.core.data_bus_o\[30\] _05028_ vssd1 vssd1 vccd1 vccd1
+ _05037_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10755__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06456__B1 total_design.core.ctrl.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_82_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12517_ net976 total_design.core.instr_mem.instruction_i\[22\] vssd1 vssd1 vccd1
+ vccd1 _01713_ sky130_fd_sc_hd__and2b_1
XANTENNA__10247__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13497_ clknet_leaf_195_clk _00964_ net1010 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12448_ net1999 net215 net344 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10771__A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09608__Y _04837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12462__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12379_ total_design.core.math.pc_val\[26\] total_design.core.program_count.imm_val_reg\[22\]
+ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07956__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11752__B2 total_design.core.data_bus_o\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14118_ clknet_leaf_101_clk _01298_ net1236 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11586__B _05479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06940_ net752 _02492_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[7\]
+ sky130_fd_sc_hd__nor2_1
X_14049_ clknet_leaf_94_clk _01229_ net1256 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11504__A1 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07708__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09771__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06399__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06871_ total_design.core.regFile.register\[3\]\[6\] net868 net761 total_design.core.regFile.register\[21\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08610_ total_design.data_in_BUS\[31\] net340 net715 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[31\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__10710__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09590_ total_design.core.ctrl.instruction\[24\] net886 net754 total_design.core.data_cpu_o\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08541_ _03875_ _03888_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08133__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09330__C1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08472_ _03798_ _03824_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07423_ total_design.core.ctrl.instruction\[29\] net887 net550 _02947_ vssd1 vssd1
+ vccd1 vccd1 _02948_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_147_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11541__S net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout147_A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07354_ total_design.core.regFile.register\[23\]\[15\] net812 net808 total_design.core.regFile.register\[5\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__a22o_1
XANTENNA__07239__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06305_ _01869_ _01882_ _01871_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12672__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10157__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07285_ total_design.core.regFile.register\[0\]\[14\] net683 _02811_ _02817_ vssd1
+ vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__o22a_2
XFILLER_0_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ net313 _04261_ _04276_ _04098_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__o211a_1
X_06236_ total_design.core.instr_mem.instruction_adr_i\[21\] total_design.core.instr_mem.instruction_adr_stored\[21\]
+ net981 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__mux2_1
XANTENNA__09946__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 total_design.lcd_display.row_1\[68\] vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
X_06167_ total_design.core.data_mem.state\[0\] vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_76_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold231 total_design.lcd_display.row_1\[91\] vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold242 total_design.lcd_display.row_1\[110\] vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold253 total_design.lcd_display.row_1\[64\] vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07947__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11743__B2 total_design.core.data_bus_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold264 total_design.lcd_display.row_1\[59\] vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07411__A2 total_design.core.data_mem.data_cpu_i\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold275 total_design.lcd_display.row_1\[3\] vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout700 _05029_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_2
Xhold286 total_design.lcd_display.row_1\[38\] vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout683_A _02035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold297 total_design.lcd_display.row_1\[117\] vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 net713 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13807__RESET_B net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout722 _02150_ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__dlymetal6s2s_1
X_09926_ net262 net2788 net424 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_165_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout733 _02037_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_2
Xfanout744 net748 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_2
Xfanout755 net756 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout766 _01997_ vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout850_A _01951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09857_ net265 net2710 net433 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__mux2_1
Xfanout777 _01990_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_8
Xfanout788 net789 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_4
XFILLER_0_137_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout799 net801 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout569_X net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10620__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ _04058_ _04060_ _04062_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__nand3_1
X_09788_ net267 net2506 net438 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__mux2_1
X_08739_ _03090_ _03138_ _03187_ _03994_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__and4_1
XANTENNA__08124__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07478__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11750_ net2876 net960 net293 total_design.core.data_bus_o\[22\] vssd1 vssd1 vccd1
+ vccd1 _01378_ sky130_fd_sc_hd__a22o_1
XANTENNA__06893__X _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10701_ net250 net2300 net359 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__mux2_1
X_11681_ _05633_ net1782 net131 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout903_X net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11451__S net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13420_ clknet_leaf_169_clk _00887_ net1160 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10632_ net275 net2580 net478 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10563_ net270 net2560 net369 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10067__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13351_ clknet_leaf_174_clk _00818_ net1054 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12302_ total_design.core.math.pc_val\[18\] total_design.core.program_count.imm_val_reg\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__and2_1
XANTENNA__09856__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06491__D net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07650__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13282_ clknet_leaf_131_clk _00749_ net1197 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10494_ net286 net2495 net481 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12233_ _06068_ _06069_ _06070_ _06076_ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11734__B2 total_design.core.data_bus_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ net1266 _01766_ _06016_ _05759_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__a31oi_1
XANTENNA__07402__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11115_ _05360_ _05368_ _05369_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_9_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12095_ total_design.lcd_display.row_1\[37\] _05827_ _05839_ total_design.lcd_display.row_1\[61\]
+ _03928_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11046_ _05295_ _05304_ _05243_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__o21bai_2
XTAP_TAPCELL_ROW_30_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11626__S net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09604__B net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10530__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08115__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08779__A_N _02718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12997_ clknet_leaf_117_clk _00464_ net1212 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11948_ _05807_ _05809_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__nor2_4
XFILLER_0_157_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06677__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12457__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11879_ net995 net897 vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__and2_2
X_13618_ clknet_leaf_48_clk net1324 net1098 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13549_ clknet_leaf_4_clk _01016_ net1022 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09766__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07070_ total_design.core.regFile.register\[26\]\[10\] net869 net846 total_design.core.regFile.register\[15\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__a22o_1
XANTENNA__07641__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10705__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07929__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06601__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07972_ total_design.core.regFile.register\[2\]\[28\] net785 net768 total_design.core.regFile.register\[7\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_71_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09711_ net704 _04934_ _04930_ _04105_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__o211a_1
X_06923_ total_design.core.regFile.register\[28\]\[7\] _01949_ net764 total_design.core.regFile.register\[6\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__a22o_1
XANTENNA__11536__S net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09642_ _03396_ _03415_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__and2b_1
XANTENNA__10440__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09514__B net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06854_ _02404_ _02406_ _02408_ _02410_ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_160_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07315__A total_design.core.ctrl.instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09573_ total_design.core.data_cpu_o\[23\] net755 _04798_ _04803_ vssd1 vssd1 vccd1
+ vccd1 _04804_ sky130_fd_sc_hd__a211o_2
X_06785_ total_design.core.ctrl.instruction\[17\] net886 vssd1 vssd1 vccd1 vccd1 _02346_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08524_ _01758_ _03843_ net932 vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11661__A0 _05663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07969__B _03467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ net933 _03782_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout431_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1173_A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07406_ total_design.core.regFile.register\[17\]\[16\] net821 net804 total_design.core.regFile.register\[8\]\[16\]
+ _02932_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__a221o_1
X_08386_ net933 _03742_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07880__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06592__C net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07337_ total_design.core.regFile.register\[8\]\[15\] net595 _02860_ _02865_ _02866_
+ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1059_X net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07268_ total_design.core.regFile.register\[10\]\[14\] net619 net611 total_design.core.regFile.register\[18\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__a22o_1
XANTENNA__07632__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06219_ total_design.core.data_adr_o\[12\] _01797_ net963 vssd1 vssd1 vccd1 vccd1
+ _01798_ sky130_fd_sc_hd__mux2_1
X_09007_ net323 _04259_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_167_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10615__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07199_ _02721_ _02723_ _02737_ net873 total_design.core.regFile.register\[0\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[12\] sky130_fd_sc_hd__o32a_4
XTAP_TAPCELL_ROW_167_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07209__B _02746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout530 _05787_ vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_2
Xfanout541 _03676_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_2
X_09909_ net185 net2128 net427 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__mux2_1
Xfanout552 net555 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_4
Xfanout563 net564 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_8
Xfanout574 net576 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11446__S net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout585 net588 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10350__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ clknet_leaf_135_clk _00387_ net1186 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout596 _02080_ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__buf_4
XANTENNA__07699__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12851_ clknet_leaf_182_clk _00318_ net1041 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11802_ net1871 _03910_ _05703_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__o21a_1
X_12782_ clknet_leaf_186_clk _00249_ net1031 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14521_ net1293 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_0_166_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06659__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11733_ net1753 net957 net290 total_design.core.data_bus_o\[5\] vssd1 vssd1 vccd1
+ vccd1 _01361_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14452_ clknet_leaf_54_clk net1351 net1110 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06275__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11664_ _05670_ net1755 net130 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13403_ clknet_leaf_143_clk _00870_ net1173 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10615_ net197 net2211 net366 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14383_ clknet_leaf_146_clk _01524_ net1178 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11595_ _05663_ net1806 net138 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07084__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13334_ clknet_leaf_155_clk _00801_ net1139 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10546_ net209 net2862 net375 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ clknet_leaf_147_clk _00732_ net1148 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10525__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10477_ net220 net2464 net379 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12216_ _06051_ _06056_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13196_ clknet_leaf_167_clk _00663_ net1155 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12147_ total_design.lcd_display.row_1\[71\] _05804_ _05810_ total_design.lcd_display.row_1\[103\]
+ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12078_ total_design.lcd_display.row_1\[76\] _05816_ _05827_ total_design.lcd_display.row_1\[36\]
+ _05935_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09533__C1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11029_ _05056_ _05275_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__and2_1
XANTENNA__10260__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06898__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11880__A total_design.core.math.pc_val\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06570_ total_design.core.regFile.register\[17\]\[1\] net822 net783 total_design.core.regFile.register\[2\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11643__A0 _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09350__A _02770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08240_ net1480 net542 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[23\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_28_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07862__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08171_ net892 _02845_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[14\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_136_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07122_ total_design.core.regFile.register\[15\]\[11\] net604 _02663_ net689 vssd1
+ vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__a211o_1
XFILLER_0_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07075__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07614__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07053_ _02596_ _02597_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06822__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10435__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07955_ _03447_ _03449_ _03451_ _03453_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__or4_1
XANTENNA__13692__D net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout381_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06906_ total_design.core.regFile.register\[15\]\[7\] net607 net582 total_design.core.regFile.register\[6\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__a22o_1
XANTENNA__10170__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07886_ total_design.core.regFile.register\[12\]\[26\] net774 net772 total_design.core.regFile.register\[28\]\[26\]
+ _03387_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__a221o_1
XANTENNA__06587__C net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07045__A total_design.core.ctrl.instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__06889__B1 total_design.core.ctrl.instruction\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_97_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09625_ _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__inv_2
X_06837_ net752 _02395_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[5\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout646_A _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09556_ _03279_ _04786_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__xor2_1
X_06768_ total_design.core.regFile.register\[20\]\[4\] net670 net593 total_design.core.regFile.register\[8\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08507_ _03837_ _03839_ _03857_ _03858_ _03768_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__o311a_1
XANTENNA__11634__A0 _05655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09487_ net211 net2602 net455 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06699_ total_design.core.ctrl.instruction\[10\] _01918_ net886 total_design.core.ctrl.instruction\[15\]
+ _02264_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__a221o_1
X_08438_ _03745_ _03765_ _03764_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_156_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07853__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08369_ total_design.keypad0.key_out\[2\] total_design.keypad0.key_out\[5\] vssd1
+ vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10400_ net259 net2302 net386 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__mux2_1
X_11380_ _05612_ _05613_ _05622_ _05638_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__and4_1
XFILLER_0_150_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07605__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13867__D total_design.core.ctrl.imm_32\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10331_ net279 net2268 net489 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__mux2_1
XANTENNA__06813__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10345__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09419__B _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13050_ clknet_leaf_125_clk _00517_ net1188 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10262_ _04112_ _04113_ _05002_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__or3_4
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout970_X net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ total_design.lcd_display.row_1\[112\] _05814_ _05838_ total_design.lcd_display.row_1\[24\]
+ _05858_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__a221o_1
XANTENNA__08030__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ _04401_ net2789 net392 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__mux2_1
Xfanout360 _05017_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_4
Xfanout371 _05013_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_6
XANTENNA__10080__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout382 net384 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_8
X_13952_ clknet_leaf_98_clk _01132_ net1242 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10125__A0 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout393 _04993_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_4
X_12903_ clknet_leaf_176_clk _00370_ net1052 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13883_ clknet_leaf_39_clk total_design.core.ctrl.imm_32\[22\] net1095 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[22\] sky130_fd_sc_hd__dfrtp_1
X_12834_ clknet_leaf_131_clk _00301_ net1197 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12704__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11625__A0 _05626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09294__A1 _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08097__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12765_ clknet_leaf_9_clk _00232_ net1020 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14504_ clknet_leaf_46_clk _01571_ vssd1 vssd1 vccd1 vccd1 total_design.key_data
+ sky130_fd_sc_hd__dfxtp_1
X_11716_ net21 net934 net877 net1635 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07844__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12696_ clknet_leaf_133_clk _00163_ net1195 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14435_ clknet_leaf_34_clk total_design.core.data_out_INSTR\[30\] net1067 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[30\] sky130_fd_sc_hd__dfrtp_1
X_11647_ _05646_ net1650 net134 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput35 gpio_in[30] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__dlymetal6s2s_1
X_14366_ clknet_leaf_122_clk _01507_ net1168 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11578_ _05648_ net1649 net142 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold808 total_design.core.regFile.register\[8\]\[3\] vssd1 vssd1 vccd1 vccd1 net2124
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06804__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13317_ clknet_leaf_117_clk _00784_ net1161 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10529_ net278 net2586 net373 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__mux2_1
XANTENNA__10255__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold819 total_design.core.regFile.register\[16\]\[6\] vssd1 vssd1 vccd1 vccd1 net2135
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_172_Right_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14297_ clknet_leaf_103_clk _00011_ net1238 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13248_ clknet_leaf_201_clk _00715_ net1004 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13179_ clknet_leaf_145_clk _00646_ net1177 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08021__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09345__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06321__X _01900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1508 total_design.core.regFile.register\[14\]\[15\] vssd1 vssd1 vccd1 vccd1 net2824
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08309__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_194_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1519 total_design.core.regFile.register\[14\]\[0\] vssd1 vssd1 vccd1 vccd1 net2835
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07740_ total_design.core.regFile.register\[10\]\[23\] net834 net775 total_design.core.regFile.register\[22\]\[23\]
+ _03236_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_88_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07671_ _03181_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__inv_2
XANTENNA__10778__X _05037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ _04128_ _04194_ _04647_ _02337_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__a22o_1
X_06622_ total_design.core.regFile.register\[30\]\[2\] net838 vssd1 vssd1 vccd1 vccd1
+ _02192_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11616__A0 _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09341_ _04571_ _04581_ net449 vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a21o_1
X_06553_ total_design.core.regFile.register\[11\]\[1\] net920 net913 net911 vssd1
+ vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_138_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08088__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09272_ total_design.core.math.pc_val\[9\] total_design.core.math.pc_val\[10\] _04471_
+ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06484_ net745 net736 net733 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__and3_1
XANTENNA__07835__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_132_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08223_ net1370 net545 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[6\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12041__B1 _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ net305 _03643_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_151_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07105_ _02637_ _02639_ _02634_ vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__o21a_1
XANTENNA__10165__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08085_ total_design.core.regFile.register\[23\]\[30\] net680 net572 total_design.core.regFile.register\[17\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_147_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1136_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09954__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07036_ total_design.core.regFile.register\[0\]\[9\] net876 _02571_ _02583_ vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[9\] sky130_fd_sc_hd__o22a_4
XFILLER_0_140_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07220__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout763_A _01997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ net469 _02367_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__nor2_1
XANTENNA__06574__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ total_design.core.regFile.register\[21\]\[27\] net761 _03434_ _03437_ vssd1
+ vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_127_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07869_ _03369_ _03370_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout551_X net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ _04827_ _04836_ net450 vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_27_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10880_ _05132_ _05138_ _05129_ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__a21o_2
XANTENNA__11607__A0 _05636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09539_ net314 _04770_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__nor2_1
XANTENNA__08079__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout816_X net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_159_Left_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12550_ net1451 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07287__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ net1586 _05679_ net151 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12481_ net982 total_design.core.instr_mem.instruction_i\[4\] vssd1 vssd1 vccd1 vccd1
+ _01695_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14220_ clknet_leaf_59_clk _01400_ net1126 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dfrtp_1
X_11432_ net1524 _05632_ net159 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__mux2_1
XANTENNA__12032__B1 _05829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09579__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ clknet_leaf_35_clk _01331_ net1068 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11363_ _05618_ _05621_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__and2_1
XANTENNA__10075__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10594__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13102_ clknet_leaf_188_clk _00569_ net1028 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09864__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10314_ net216 net2675 net492 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__mux2_1
X_14082_ clknet_leaf_87_clk _01262_ net1248 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[36\]
+ sky130_fd_sc_hd__dfrtp_1
X_11294_ _05545_ _05546_ _05551_ _05515_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__o22ai_2
XPHY_EDGE_ROW_168_Left_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08988__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13033_ clknet_leaf_19_clk _00500_ net1050 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08003__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10245_ net226 net2473 net502 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__mux2_1
Xfanout1100 net1104 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1111 net1121 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__clkbuf_4
Xfanout1122 net1123 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__clkbuf_4
X_10176_ net203 net1954 net395 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__mux2_1
Xfanout1133 net1134 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__clkbuf_2
Xfanout1144 net1172 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__buf_2
XANTENNA__06565__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1155 net1163 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12099__B1 _05838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1166 net1168 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__clkbuf_4
Xfanout1177 net1178 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__clkbuf_4
Xfanout190 net192 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_1
Xfanout1188 net1190 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__clkbuf_4
Xfanout1199 net1200 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__clkbuf_2
X_13935_ clknet_leaf_84_clk _01115_ net1245 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11634__S net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13866_ clknet_leaf_65_clk total_design.core.ctrl.imm_32\[5\] net1124 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12817_ clknet_leaf_152_clk _00284_ net1146 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13797_ clknet_4_13__leaf_clk total_design.core.data_mem.data_cpu_i\[6\] net1212
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08228__B net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11074__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12748_ clknet_leaf_165_clk _00215_ net1157 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10774__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12679_ clknet_leaf_173_clk _00146_ net1052 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14418_ clknet_leaf_36_clk total_design.core.data_out_INSTR\[13\] net1071 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[13\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12023__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14349_ clknet_leaf_45_clk _00036_ net1088 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold605 total_design.core.regFile.register\[25\]\[6\] vssd1 vssd1 vccd1 vccd1 net1921
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 total_design.core.regFile.register\[19\]\[19\] vssd1 vssd1 vccd1 vccd1 net1932
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09774__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold627 total_design.core.regFile.register\[31\]\[12\] vssd1 vssd1 vccd1 vccd1 net1943
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 total_design.core.regFile.register\[17\]\[21\] vssd1 vssd1 vccd1 vccd1 net1954
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07450__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold649 total_design.core.regFile.register\[18\]\[13\] vssd1 vssd1 vccd1 vccd1 net1965
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08910_ net471 net305 _04163_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12053__X _05912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10713__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09890_ net274 net1921 net428 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08841_ _04086_ _04089_ _04095_ _04074_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__o31a_1
Xhold1305 total_design.core.regFile.register\[11\]\[18\] vssd1 vssd1 vccd1 vccd1 net2621
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1316 total_design.core.regFile.register\[27\]\[7\] vssd1 vssd1 vccd1 vccd1 net2632
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1327 total_design.core.regFile.register\[19\]\[3\] vssd1 vssd1 vccd1 vccd1 net2643
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07307__B _02818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08772_ _03486_ _03506_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__nand2_1
Xhold1338 total_design.core.regFile.register\[25\]\[2\] vssd1 vssd1 vccd1 vccd1 net2654
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1349 total_design.core.regFile.register\[27\]\[30\] vssd1 vssd1 vccd1 vccd1 net2665
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07723_ _03093_ _03136_ _03231_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11544__S net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07654_ total_design.core.regFile.register\[9\]\[21\] net664 net621 total_design.core.regFile.register\[4\]\[21\]
+ _03164_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06605_ total_design.core.regFile.register\[27\]\[1\] net580 _02157_ _02161_ _02164_
+ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_88_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07585_ total_design.core.regFile.register\[29\]\[20\] net655 net566 total_design.core.regFile.register\[12\]\[20\]
+ _03098_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout344_A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1086_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09949__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06584__D net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07269__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ _02718_ _02738_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__nand2_1
X_06536_ total_design.core.ctrl.imm_32\[0\] _02109_ vssd1 vssd1 vccd1 vccd1 _02110_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07808__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08853__S _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09255_ _02637_ _04498_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout132_X net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout511_A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06467_ total_design.core.regFile.register\[22\]\[0\] net747 net735 net731 vssd1
+ vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__and4_1
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout609_A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ _03659_ _03660_ _03662_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__or3_1
XFILLER_0_145_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13414__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12014__B1 _05840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06398_ net922 net919 net914 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__and3_1
X_09186_ _04322_ _04324_ net329 vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08154__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08137_ total_design.core.regFile.register\[24\]\[31\] net574 net571 total_design.core.regFile.register\[17\]\[31\]
+ _03624_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07441__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08068_ total_design.core.regFile.register\[10\]\[30\] net836 net792 total_design.core.regFile.register\[24\]\[30\]
+ _03561_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout978_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06795__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07019_ total_design.core.regFile.register\[30\]\[9\] net840 net778 total_design.core.regFile.register\[22\]\[9\]
+ _02566_ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__a221o_1
XANTENNA__10623__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ net255 net2535 net410 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06402__A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11962__B _05823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ _05754_ _05842_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__nor2_4
XANTENNA__13880__D total_design.core.ctrl.imm_32\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13720_ clknet_leaf_35_clk total_design.core.data_mem.stored_read_data\[27\] net1068
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[27\] sky130_fd_sc_hd__dfrtp_1
X_10932_ _05183_ _05188_ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13651_ clknet_leaf_50_clk total_design.core.data_mem.data_write_adr_i\[23\] net1100
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[23\] sky130_fd_sc_hd__dfrtp_1
X_10863_ _05099_ _05101_ _05102_ vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12602_ clknet_leaf_125_clk _00069_ net1189 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09859__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13582_ clknet_leaf_34_clk total_design.core.data_mem.data_bus_i\[18\] net1066 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[18\] sky130_fd_sc_hd__dfrtp_1
X_10794_ _05049_ _05052_ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12533_ net974 total_design.core.instr_mem.instruction_i\[30\] vssd1 vssd1 vccd1
+ vccd1 _01721_ sky130_fd_sc_hd__and2b_1
XFILLER_0_109_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12005__B1 _05830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06283__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12464_ _03985_ _05784_ total_design.keypad0.key_counter\[0\] vssd1 vssd1 vccd1 vccd1
+ _01686_ sky130_fd_sc_hd__o21a_1
XANTENNA__07680__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14203_ clknet_leaf_80_clk _01383_ net1222 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
X_11415_ _05609_ _05639_ _05649_ _05673_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__and4_2
XFILLER_0_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12395_ net899 _03467_ net523 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14134_ clknet_leaf_101_clk _01314_ net1240 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07432__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11346_ _05450_ _05452_ _05454_ _05465_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11629__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14065_ clknet_leaf_94_clk _01245_ net1256 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10533__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09166__Y _04414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ _05442_ _05447_ _05535_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__nand3_1
X_13016_ clknet_leaf_146_clk _00483_ net1178 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10228_ total_design.core.ctrl.instruction\[11\] net556 total_design.core.instr_fetch
+ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_33_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 total_design.core.instr_mem.instr_fetch vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ net280 net2829 net394 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07499__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13918_ clknet_leaf_96_clk _01098_ net1254 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13849_ clknet_leaf_48_clk _01057_ net1099 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06710__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09769__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07370_ net550 _02896_ _02897_ vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[16\]
+ sky130_fd_sc_hd__or3b_2
XFILLER_0_57_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06321_ _01891_ _01893_ _01898_ _01899_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__and4_2
XFILLER_0_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10708__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06252_ total_design.core.instr_mem.instruction_adr_i\[22\] total_design.core.instr_mem.instruction_adr_stored\[22\]
+ net981 vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__mux2_1
X_09040_ net535 _04285_ _04291_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06183_ total_design.bus_full _01730_ total_design.key_data vssd1 vssd1 vccd1 vccd1
+ _01764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold402 total_design.lcd_display.row_2\[32\] vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 total_design.lcd_display.row_2\[46\] vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold424 net44 vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold435 total_design.lcd_display.row_1\[79\] vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 total_design.lcd_display.row_2\[87\] vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold457 total_design.lcd_display.row_2\[13\] vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 total_design.lcd_display.row_2\[104\] vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09942_ net189 net2272 net423 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold479 net41 vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10443__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout904 net905 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__buf_4
Xfanout915 _01937_ vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_74_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout926 _01925_ vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_2
Xfanout937 _05688_ vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__dlymetal6s2s_1
X_09873_ net196 net2009 net430 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__mux2_1
Xfanout948 _01929_ vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__buf_2
XANTENNA__06529__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 net960 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 total_design.core.regFile.register\[13\]\[22\] vssd1 vssd1 vccd1 vccd1 net2418
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08824_ _04072_ _04077_ _04078_ _04057_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__a31o_1
Xhold1113 total_design.core.regFile.register\[21\]\[19\] vssd1 vssd1 vccd1 vccd1 net2429
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1124 total_design.core.regFile.register\[12\]\[22\] vssd1 vssd1 vccd1 vccd1 net2440
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1135 total_design.core.regFile.register\[5\]\[21\] vssd1 vssd1 vccd1 vccd1 net2451
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 total_design.core.regFile.register\[20\]\[22\] vssd1 vssd1 vccd1 vccd1 net2462
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1157 total_design.core.regFile.register\[15\]\[15\] vssd1 vssd1 vccd1 vccd1 net2473
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ _02968_ net309 _04008_ _04009_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__a211o_1
Xhold1168 total_design.core.regFile.register\[21\]\[14\] vssd1 vssd1 vccd1 vccd1 net2484
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 total_design.core.regFile.register\[7\]\[0\] vssd1 vssd1 vccd1 vccd1 net2495
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ total_design.core.regFile.register\[25\]\[22\] net648 net586 total_design.core.regFile.register\[28\]\[22\]
+ _03210_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__a221o_1
X_08686_ _03960_ _03961_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06595__C net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07637_ total_design.core.regFile.register\[18\]\[21\] net859 _03146_ _03147_ _03148_
+ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_95_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout726_A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07568_ _03064_ _03084_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__nand2_1
XANTENNA__06892__A total_design.core.ctrl.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09307_ _04132_ _04137_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__or2_1
X_06519_ total_design.core.regFile.register\[12\]\[0\] _02031_ net739 net727 vssd1
+ vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__and4_1
XFILLER_0_1_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10618__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07499_ total_design.core.regFile.register\[31\]\[18\] net831 net806 total_design.core.regFile.register\[5\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08155__Y _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07662__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09238_ _04439_ _04482_ net463 vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10549__A0 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09403__A1 _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ _04416_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11200_ net303 vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__inv_2
X_12180_ _06029_ _06030_ net994 vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06768__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11449__S net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11761__A2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ _05386_ _05388_ _05380_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_102_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10353__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 total_design.core.regFile.register\[7\]\[14\] vssd1 vssd1 vccd1 vccd1 net2296
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 total_design.core.regFile.register\[1\]\[24\] vssd1 vssd1 vccd1 vccd1 net2307
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ net352 _05063_ _05264_ _05314_ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__a2bb2o_1
X_10013_ net176 net2678 net417 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__mux2_1
XANTENNA__06489__D net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07193__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06278__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12474__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11964_ _05811_ _05825_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__nor2_4
XANTENNA__08059__A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13703_ clknet_leaf_38_clk total_design.core.data_mem.stored_read_data\[10\] net1079
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[10\] sky130_fd_sc_hd__dfrtp_1
X_10915_ _05172_ _05173_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11895_ net35 net38 net37 net36 vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__or4b_1
XFILLER_0_129_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13634_ clknet_leaf_60_clk total_design.core.data_mem.data_write_adr_i\[6\] net1131
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10846_ _05099_ _05104_ _05089_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13565_ clknet_leaf_38_clk total_design.core.data_mem.data_bus_i\[1\] net1078 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[1\] sky130_fd_sc_hd__dfrtp_1
X_10777_ total_design.core.data_bus_o\[19\] net695 vssd1 vssd1 vccd1 vccd1 _05036_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10528__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12516_ net976 total_design.core.ctrl.instruction\[21\] net881 _01712_ vssd1 vssd1
+ vccd1 vccd1 _01560_ sky130_fd_sc_hd__a22o_1
XANTENNA__07653__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06307__A _01852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13496_ clknet_leaf_135_clk _00963_ net1189 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12447_ net1883 net220 net346 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__mux2_1
XANTENNA__09177__X _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07405__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12378_ total_design.core.math.pc_val\[26\] total_design.core.program_count.imm_val_reg\[22\]
+ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06759__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14117_ clknet_leaf_88_clk _01297_ net1251 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11329_ _05578_ _05584_ _05586_ _05587_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__or4_1
XANTENNA__10263__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09158__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14048_ clknet_leaf_110_clk _01228_ net1227 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06870_ total_design.core.regFile.register\[16\]\[6\] net856 net785 total_design.core.regFile.register\[2\]\[6\]
+ _02426_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07184__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06931__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08540_ _03875_ _03888_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08471_ _03823_ _03801_ net931 vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07422_ _02945_ _02946_ net721 vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07353_ total_design.core.regFile.register\[12\]\[15\] net774 net772 total_design.core.regFile.register\[28\]\[15\]
+ _02882_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__a221o_1
XANTENNA__10438__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06304_ _01869_ _01882_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__and2_1
XANTENNA__11440__A1 _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07284_ _02813_ _02814_ _02815_ _02816_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__or4_1
XFILLER_0_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06998__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14207__Q net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09023_ net313 _04275_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__nand2_1
X_06235_ net929 _01813_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10962__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1049_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 total_design.lcd_display.row_1\[12\] vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_1__f_clk_X clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06166_ net1626 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__inv_2
Xhold221 total_design.lcd_display.row_1\[0\] vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold232 total_design.lcd_display.row_1\[113\] vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold243 net69 vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11743__A2 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold254 total_design.lcd_display.row_1\[39\] vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10173__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold265 total_design.lcd_display.row_1\[15\] vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold276 total_design.core.math.pc_val\[21\] vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold287 total_design.lcd_display.row_1\[33\] vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout701 net702 vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__buf_2
XANTENNA__09962__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold298 total_design.lcd_display.row_2\[116\] vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ net266 net1996 net422 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__mux2_1
XANTENNA__09815__X _04973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout712 net713 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_1
Xfanout723 net725 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout734 net735 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_123_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout676_A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 net748 vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_1
XANTENNA_fanout297_X net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout756 net757 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout767 net770 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__buf_4
X_09856_ net273 net2443 net431 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1004_X net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout778 _01990_ vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06887__A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout789 _01984_ vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_4
X_08807_ _04059_ _04061_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__and2b_1
X_09787_ net272 net2521 net440 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout843_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06999_ total_design.core.regFile.register\[15\]\[9\] net606 net584 total_design.core.regFile.register\[6\]\[9\]
+ _02546_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a221o_1
XANTENNA__06922__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ _02944_ _02993_ _03040_ _03993_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__and4_1
XFILLER_0_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09550__X _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08669_ total_design.lcd_display.cnt_500hz\[13\] _03946_ _03947_ vssd1 vssd1 vccd1
+ vccd1 _00009_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout729_X net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10700_ net261 net2252 net360 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__mux2_1
X_11680_ _05646_ net1841 net130 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__mux2_1
XANTENNA__07883__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10631_ net259 net2156 net478 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10348__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11431__A1 _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07635__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ clknet_leaf_197_clk _00817_ net1007 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10562_ net277 net2026 net369 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12301_ total_design.core.math.pc_val\[17\] net524 _06137_ _06138_ vssd1 vssd1 vccd1
+ vccd1 _01487_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13281_ clknet_leaf_123_clk _00748_ net1167 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10493_ _04972_ _04980_ _05002_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__or3_4
XFILLER_0_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12232_ _06068_ _06069_ _06070_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_20_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06414__X _01990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12163_ total_design.core.disable_pc_reg total_design.core.data_access vssd1 vssd1
+ vccd1 vccd1 _06016_ sky130_fd_sc_hd__nor2_1
XANTENNA__10083__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09872__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ _05368_ _05369_ _05360_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_9_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09725__X _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12094_ total_design.lcd_display.row_2\[85\] _05818_ _05853_ total_design.lcd_display.row_2\[117\]
+ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__a22o_1
X_11045_ _05056_ _05299_ _05300_ _05303_ _05298_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11498__A1 _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07166__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06374__B1 total_design.core.ctrl.instruction\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12996_ clknet_leaf_106_clk _00463_ net1223 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_12__f_clk_X clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11947_ _05754_ _05808_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__or2_4
XFILLER_0_8_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11642__S net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07874__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ total_design.core.disable_pc_reg _05757_ vssd1 vssd1 vccd1 vccd1 _05759_
+ sky130_fd_sc_hd__nor2_1
X_13617_ clknet_leaf_47_clk net1346 net1098 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10829_ _05061_ _05086_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__nor2_1
XANTENNA__10258__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13548_ clknet_leaf_169_clk _01015_ net1160 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13479_ clknet_leaf_177_clk _00946_ net1047 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14549__1269 vssd1 vssd1 vccd1 vccd1 _14549__1269/HI net1269 sky130_fd_sc_hd__conb_1
XANTENNA__09348__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09782__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07971_ total_design.core.regFile.register\[12\]\[28\] net773 net771 total_design.core.regFile.register\[28\]\[28\]
+ _03468_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_71_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09710_ _03600_ _04932_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_143_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06922_ total_design.core.regFile.register\[1\]\[7\] net827 net759 total_design.core.regFile.register\[21\]\[7\]
+ _02475_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_143_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10721__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12150__A2 _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ _03467_ net707 vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__or2_1
XANTENNA__07011__D1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06853_ total_design.core.regFile.register\[19\]\[6\] net642 net614 total_design.core.regFile.register\[11\]\[6\]
+ _02409_ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_160_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06904__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09572_ net965 net886 _04802_ net906 vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__a22o_1
X_06784_ total_design.core.ctrl.instruction\[25\] _02312_ vssd1 vssd1 vccd1 vccd1
+ _02345_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08523_ net717 _03873_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[9\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_69_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11552__S net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06668__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ net933 total_design.keypad0.key_out\[8\] vssd1 vssd1 vccd1 vccd1 _03808_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_0_147_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07405_ total_design.core.regFile.register\[26\]\[16\] net871 net848 total_design.core.regFile.register\[15\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__a22o_1
X_08385_ _03739_ _03740_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__xor2_1
XANTENNA__10168__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout424_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09957__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ total_design.core.regFile.register\[7\]\[15\] net654 net642 total_design.core.regFile.register\[19\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07267_ total_design.core.regFile.register\[30\]\[14\] net662 _02076_ total_design.core.regFile.register\[31\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_115_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09006_ _04255_ _04258_ net468 vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06218_ total_design.core.instr_mem.instruction_adr_i\[12\] total_design.core.instr_mem.instruction_adr_stored\[12\]
+ net983 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07198_ _02726_ _02728_ _02730_ _02736_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_167_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06149_ total_design.keypad0.key_out\[3\] vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08042__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1121_X net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07396__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout960_A _01911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout581_X net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout520 _01885_ vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_4
Xfanout531 _05755_ vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout542 net544 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_2
X_09908_ net191 net2751 net428 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__mux2_1
XANTENNA__10631__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout553 net554 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_4
Xfanout564 net565 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__buf_4
Xfanout575 net576 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_4
XANTENNA__12141__A2 _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout586 net588 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_8
X_09839_ net195 net2118 net434 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__mux2_1
Xfanout597 net600 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06410__A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout846_X net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ clknet_leaf_139_clk _00317_ net1184 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11801_ _03912_ net713 vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12781_ clknet_leaf_0_clk _00248_ net1004 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11462__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_140_Left_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14520_ net1292 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
X_11732_ net1843 net957 net290 total_design.core.data_bus_o\[4\] vssd1 vssd1 vccd1
+ vccd1 _01360_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07856__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07320__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14451_ clknet_leaf_67_clk net1731 net1122 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11663_ _05667_ net1730 net129 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__mux2_1
XANTENNA__10078__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09058__C1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ clknet_leaf_132_clk _00869_ net1196 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10614_ net203 net2045 net366 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__mux2_1
XANTENNA__07608__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09867__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14382_ clknet_leaf_150_clk _01523_ net1147 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11594_ _05627_ net1654 net140 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13333_ clknet_leaf_160_clk _00800_ net1142 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10545_ net217 net2590 net373 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_130_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13264_ clknet_leaf_185_clk _00731_ net1038 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10476_ net226 net2338 net379 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12215_ _06060_ _06061_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__nand2_1
XANTENNA__08033__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13195_ clknet_leaf_107_clk _00662_ net1224 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07387__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09455__X _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ total_design.lcd_display.row_1\[127\] _05843_ _05853_ total_design.lcd_display.row_2\[119\]
+ _06000_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__a221o_1
XANTENNA__11637__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10541__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12077_ total_design.lcd_display.row_1\[84\] _05815_ _05932_ _05934_ vssd1 vssd1
+ vccd1 vccd1 _05935_ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07139__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11028_ _05274_ _05277_ _05269_ _05270_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__o211ai_2
XANTENNA__06320__A _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_197_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_197_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06347__B1 _01915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12979_ clknet_leaf_179_clk _00446_ net1035 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09777__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ net892 _02796_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[13\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_136_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07121_ total_design.core.regFile.register\[11\]\[11\] net615 net585 total_design.core.regFile.register\[28\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10716__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_121_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11401__A _05651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07052_ total_design.core.regFile.register\[13\]\[10\] net666 net562 total_design.core.regFile.register\[3\]\[10\]
+ _02594_ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a221o_1
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__clkbuf_4
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_11_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__08024__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07378__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10451__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07954_ total_design.core.regFile.register\[16\]\[27\] net635 net583 total_design.core.regFile.register\[6\]\[27\]
+ _03452_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__a221o_1
XANTENNA__12123__A2 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06905_ total_design.core.regFile.register\[14\]\[7\] net627 net588 total_design.core.regFile.register\[28\]\[7\]
+ _02458_ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a221o_1
X_07885_ total_design.core.regFile.register\[20\]\[26\] net816 net815 total_design.core.regFile.register\[4\]\[26\]
+ net692 vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_188_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_188_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout374_A _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ _04166_ _04168_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__nor2_1
X_06836_ _02348_ _02394_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__xor2_2
XANTENNA__06587__D net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07550__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13021__RESET_B net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09555_ _04762_ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__or2_1
X_06767_ _02322_ _02324_ _02326_ _02328_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout541_A _03676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06884__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08506_ _03837_ _03839_ _03857_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__o21ai_1
X_09486_ net507 _04720_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__and2_1
X_06698_ net949 net947 _02149_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__o21a_1
XANTENNA__07302__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08437_ _03790_ _03791_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout806_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08368_ total_design.keypad0.key_out\[2\] total_design.keypad0.key_out\[5\] vssd1
+ vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07319_ _02839_ _02843_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__and2b_1
XANTENNA__10626__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08299_ total_design.core.data_mem.data_write_adr_reg\[7\] net549 net541 total_design.core.data_mem.data_read_adr_reg\[7\]
+ net945 vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_112_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12407__A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10330_ net246 net2877 net491 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout796_X net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ net162 net2600 net501 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12000_ _05855_ _05857_ _05860_ _05861_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__or4_1
X_10192_ net282 net1908 net389 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout963_X net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11570__A0 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11457__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout350 _05044_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_2
Xfanout361 net364 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09515__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout372 _05013_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_4
X_13951_ clknet_leaf_84_clk _01131_ net1245 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[33\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_179_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_179_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout383 net384 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout394 net397 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_6
X_12902_ clknet_leaf_200_clk _00369_ net1002 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13882_ clknet_leaf_38_clk total_design.core.ctrl.imm_32\[21\] net1079 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[21\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09451__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07541__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14548__1268 vssd1 vssd1 vccd1 vccd1 _14548__1268/HI net1268 sky130_fd_sc_hd__conb_1
X_12833_ clknet_leaf_164_clk _00300_ net1165 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07829__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12764_ clknet_leaf_29_clk _00231_ net1063 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11715_ net20 net936 net879 net1832 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__a22o_1
X_14503_ clknet_leaf_27_clk _01570_ net1077 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_139_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12695_ clknet_leaf_166_clk _00162_ net1164 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11646_ _05645_ net1638 net133 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__mux2_1
X_14434_ clknet_leaf_36_clk total_design.core.data_out_INSTR\[29\] net1072 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[29\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14365_ clknet_leaf_194_clk _01506_ net1011 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
X_11577_ _05628_ net1766 net143 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__mux2_1
Xinput36 gpio_in[31] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
XANTENNA__10536__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_103_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11221__A _05479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13316_ clknet_leaf_128_clk _00783_ net1194 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10528_ net247 net2239 net374 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__mux2_1
Xhold809 total_design.core.regFile.register\[28\]\[28\] vssd1 vssd1 vccd1 vccd1 net2125
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14296_ clknet_leaf_103_clk _00005_ net1238 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13247_ clknet_leaf_157_clk _00714_ net1140 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08006__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10459_ net164 net2421 net383 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13178_ clknet_leaf_133_clk _00645_ net1196 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11561__A0 _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13793__D total_design.core.data_mem.data_cpu_i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12129_ total_design.lcd_display.row_1\[86\] _05815_ _05816_ total_design.lcd_display.row_1\[78\]
+ _05972_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a221o_1
XANTENNA__13532__RESET_B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10271__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1509 total_design.core.regFile.register\[9\]\[0\] vssd1 vssd1 vccd1 vccd1 net2825
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12105__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09506__B1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07780__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07670_ net299 _03180_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__nor2_1
XANTENNA__09632__Y _04860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06621_ total_design.core.regFile.register\[25\]\[2\] net845 net791 total_design.core.regFile.register\[24\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__a22o_1
XANTENNA__09361__A _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06740__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09340_ _04194_ _04575_ _04577_ _04580_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__o211a_1
X_06552_ total_design.core.regFile.register\[1\]\[1\] net921 net948 net909 vssd1 vssd1
+ vccd1 vccd1 _02125_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_138_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09271_ _04502_ _04512_ _04514_ net449 vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_103_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06483_ total_design.core.regFile.register\[26\]\[0\] net748 net730 net725 vssd1
+ vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08222_ net1361 net545 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[5\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_117_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08153_ net305 _03643_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__and2_1
XANTENNA__10446__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07104_ _02646_ vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[11\] sky130_fd_sc_hd__inv_2
XFILLER_0_130_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07599__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08084_ total_design.core.regFile.register\[2\]\[30\] net638 net622 total_design.core.regFile.register\[4\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07035_ _02576_ _02578_ _02579_ _02582_ vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout1031_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1129_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout589_A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ _04237_ _04238_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__nor2_1
XANTENNA__09970__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06598__C net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07937_ total_design.core.regFile.register\[2\]\[27\] net784 _03435_ _03436_ vssd1
+ vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout756_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07868_ _03369_ _03370_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_127_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09607_ net297 _04489_ _04667_ _04485_ _04835_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__o221a_1
X_06819_ total_design.core.regFile.register\[15\]\[5\] net848 _02378_ vssd1 vssd1
+ vccd1 vccd1 _02379_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_27_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07799_ total_design.core.regFile.register\[18\]\[24\] net609 net578 total_design.core.regFile.register\[27\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__a22o_1
XANTENNA__06731__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout923_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09538_ _04692_ _04769_ net332 vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09469_ _03090_ net703 _04703_ net533 vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout809_X net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ net1604 _05632_ net150 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__mux2_1
X_12480_ net979 total_design.core.ctrl.instruction\[3\] net884 _01694_ vssd1 vssd1
+ vccd1 vccd1 _01542_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11431_ net1530 _05670_ net160 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10356__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14150_ clknet_leaf_35_clk _01330_ net1068 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11362_ _05452_ net303 _05619_ _05620_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__o22a_2
XFILLER_0_21_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06798__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13101_ clknet_leaf_5_clk _00568_ net1022 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10313_ net213 net2682 net492 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14081_ clknet_leaf_97_clk _01261_ net1246 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11293_ _05543_ _05550_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__or2_1
X_13032_ clknet_leaf_24_clk _00499_ net1108 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10244_ net233 total_design.core.regFile.register\[15\]\[14\] net503 vssd1 vssd1
+ vccd1 vccd1 _00533_ sky130_fd_sc_hd__mux2_1
Xfanout1101 net1104 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_2
Xfanout1112 net1121 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10091__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10175_ net205 net2088 net394 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__mux2_1
Xfanout1123 net1134 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__buf_2
Xfanout1134 net1135 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__buf_2
Xfanout1145 net1149 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07762__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09880__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11982__Y _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1156 net1163 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__buf_2
Xfanout1167 net1168 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__clkbuf_4
Xfanout1178 net1181 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06970__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 net192 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_2
Xfanout1189 net1190 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__clkbuf_4
X_13934_ clknet_leaf_100_clk _01114_ net1254 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07514__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07253__X total_design.core.data_mem.data_cpu_i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13865_ clknet_leaf_65_clk total_design.core.ctrl.imm_32\[4\] net1124 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06722__B1 _02266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11059__C1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12816_ clknet_leaf_182_clk _00283_ net1041 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13796_ clknet_leaf_71_clk total_design.core.data_mem.data_cpu_i\[5\] net1205 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09267__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10806__C1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11074__A2 _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12271__A1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12747_ clknet_leaf_120_clk _00214_ net1191 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11650__S net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12678_ clknet_leaf_198_clk _00145_ net1008 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10774__B total_design.core.data_bus_o\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11629_ _05665_ net1749 net135 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__mux2_1
X_14417_ clknet_leaf_36_clk total_design.core.data_out_INSTR\[12\] net1078 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10266__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08244__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14348_ clknet_leaf_46_clk _00035_ net1088 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold606 total_design.core.regFile.register\[9\]\[16\] vssd1 vssd1 vccd1 vccd1 net1922
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06789__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold617 total_design.core.regFile.register\[18\]\[25\] vssd1 vssd1 vccd1 vccd1 net1933
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11886__A total_design.core.math.pc_val\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold628 total_design.core.regFile.register\[3\]\[7\] vssd1 vssd1 vccd1 vccd1 net1944
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10790__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14279_ net986 _01455_ net1087 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[8\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold639 total_design.core.regFile.register\[13\]\[13\] vssd1 vssd1 vccd1 vccd1 net1955
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_59_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _04090_ _04094_ _04031_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_55_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07753__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1306 total_design.core.regFile.register\[3\]\[11\] vssd1 vssd1 vccd1 vccd1 net2622
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1317 total_design.core.regFile.register\[18\]\[24\] vssd1 vssd1 vccd1 vccd1 net2633
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08771_ _04024_ _04025_ _04023_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__and3b_1
Xhold1328 total_design.core.regFile.register\[31\]\[29\] vssd1 vssd1 vccd1 vccd1 net2644
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1339 total_design.core.regFile.register\[21\]\[11\] vssd1 vssd1 vccd1 vccd1 net2655
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07722_ _03134_ _03182_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07505__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ total_design.core.regFile.register\[19\]\[21\] net641 net609 total_design.core.regFile.register\[18\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06713__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06604_ total_design.core.regFile.register\[30\]\[1\] net662 _02153_ _02155_ _02169_
+ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_0_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07584_ total_design.core.regFile.register\[4\]\[20\] net620 net577 total_design.core.regFile.register\[27\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__a22o_1
XANTENNA__09258__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09323_ net238 net1973 net456 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06535_ total_design.core.data_mem.data_cpu_i\[0\] net552 vssd1 vssd1 vccd1 vccd1
+ _02109_ sky130_fd_sc_hd__and2_1
XFILLER_0_158_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11560__S net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ _02588_ _04477_ _04497_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_29_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06466_ net744 net734 net730 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__and3_1
XFILLER_0_173_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08205_ total_design.core.data_mem.data_read_adr_reg\[29\] total_design.core.data_mem.data_read_adr_reg\[28\]
+ total_design.core.data_mem.data_read_adr_reg\[31\] total_design.core.data_mem.data_read_adr_reg\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__or4_1
XFILLER_0_106_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10176__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09185_ net322 _04321_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout504_A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06397_ total_design.core.regFile.register\[5\]\[0\] net922 _01950_ net907 vssd1
+ vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_170_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1246_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08136_ total_design.core.regFile.register\[7\]\[31\] net653 net598 total_design.core.regFile.register\[21\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__a22o_1
XANTENNA__09965__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11773__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08067_ total_design.core.regFile.register\[18\]\[30\] net859 net821 total_design.core.regFile.register\[17\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07992__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07018_ total_design.core.regFile.register\[15\]\[9\] net848 net792 total_design.core.regFile.register\[24\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__a22o_1
XANTENNA__07338__X _02868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08170__A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout873_A _01934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1201_X net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ net336 _02818_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06952__B1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11980_ _05746_ _05749_ _05813_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__or3_4
XFILLER_0_98_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10931_ _05151_ _05152_ _05189_ _05157_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__o31a_1
XANTENNA__06704__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13650_ clknet_leaf_47_clk total_design.core.data_mem.data_write_adr_i\[22\] net1097
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[22\] sky130_fd_sc_hd__dfrtp_1
X_10862_ _05115_ _05117_ _05119_ _05106_ _05105_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12601_ clknet_leaf_196_clk _00068_ net1009 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12253__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13581_ clknet_leaf_32_clk total_design.core.data_mem.data_bus_i\[17\] net1062 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[17\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10875__A _01885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10793_ total_design.core.data_bus_o\[8\] total_design.core.data_bus_o\[9\] _05050_
+ _05051_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__or4b_1
XFILLER_0_67_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11470__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10264__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12532_ net977 total_design.core.ctrl.instruction\[29\] net882 _01720_ vssd1 vssd1
+ vccd1 vccd1 _01568_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07520__Y _03040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12463_ net1834 _03975_ net1087 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_193_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11414_ _05650_ _05660_ _05668_ _05672_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__and4_1
XFILLER_0_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09875__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14202_ clknet_leaf_111_clk _01382_ net1208 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_2
XANTENNA__11977__Y _05839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12394_ net992 _01651_ _01652_ _01653_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14133_ clknet_leaf_85_clk _01313_ net1258 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11345_ _05450_ _05465_ _05603_ _05455_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_1_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07983__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14064_ clknet_leaf_109_clk _01244_ net1226 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[82\]
+ sky130_fd_sc_hd__dfrtp_1
X_11276_ _05438_ _05531_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_37_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13015_ clknet_leaf_166_clk _00482_ net1164 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10227_ total_design.core.ctrl.instruction\[11\] net556 total_design.core.instr_fetch
+ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07361__A_N _02868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07735__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10158_ net270 net2057 net395 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_131_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 total_design.core.data_mem.data_read_adr_reg\[25\] vssd1 vssd1 vccd1 vccd1
+ net1319 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11645__S net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10089_ net278 net2505 net403 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13917_ clknet_leaf_89_clk _01097_ net1258 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_146_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13848_ clknet_leaf_52_clk _01056_ net1094 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wire305_A _03642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13779_ clknet_leaf_48_clk total_design.core.data_mem.stored_data_adr\[22\] net1102
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[22\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06320_ _01808_ _01830_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06251_ total_design.core.data_adr_o\[13\] net961 net929 _01829_ vssd1 vssd1 vccd1
+ vccd1 _01830_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09785__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09638__X _04866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06182_ _01762_ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__inv_2
XANTENNA__06322__C_N _01900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold403 total_design.lcd_display.row_2\[89\] vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold414 total_design.lcd_display.row_2\[10\] vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 total_design.lcd_display.row_2\[66\] vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold436 total_design.lcd_display.row_2\[64\] vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 net43 vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold458 total_design.lcd_display.row_2\[5\] vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07974__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold469 net103 vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ net194 net2642 net422 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout905 _02015_ vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout916 _01935_ vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__buf_2
Xfanout927 net928 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__buf_2
X_09872_ net199 net2606 net431 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout938 _03675_ vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__clkbuf_4
Xfanout949 _01929_ vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 total_design.core.regFile.register\[16\]\[29\] vssd1 vssd1 vccd1 vccd1 net2419
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08823_ _04064_ _04066_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__or2_1
XANTENNA__09814__A total_design.core.ctrl.instruction\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1114 total_design.core.regFile.register\[27\]\[27\] vssd1 vssd1 vccd1 vccd1 net2430
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11555__S net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1125 total_design.core.regFile.register\[26\]\[15\] vssd1 vssd1 vccd1 vccd1 net2441
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1136 total_design.core.regFile.register\[9\]\[4\] vssd1 vssd1 vccd1 vccd1 net2452
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1147 total_design.core.regFile.register\[16\]\[12\] vssd1 vssd1 vccd1 vccd1 net2463
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ _03064_ _03083_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__and2_1
Xhold1158 total_design.core.regFile.register\[5\]\[14\] vssd1 vssd1 vccd1 vccd1 net2474
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 total_design.core.regFile.register\[3\]\[4\] vssd1 vssd1 vccd1 vccd1 net2485
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ total_design.core.regFile.register\[13\]\[22\] net667 net637 total_design.core.regFile.register\[2\]\[22\]
+ _03211_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08685_ total_design.keypad0.counter\[16\] _03958_ net2612 vssd1 vssd1 vccd1 vccd1
+ _03961_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_92_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_135_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout454_A _04117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08151__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10494__A0 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07636_ total_design.core.regFile.register\[19\]\[21\] net824 net780 total_design.core.regFile.register\[27\]\[21\]
+ _03139_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_120_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12235__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07567_ net552 total_design.core.data_mem.data_cpu_i\[19\] total_design.core.ctrl.imm_32\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_172_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout621_A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09306_ net702 _04546_ _04547_ _04105_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout719_A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06518_ net740 net739 net726 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__and3_4
XANTENNA__08165__A _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07498_ total_design.core.regFile.register\[15\]\[18\] net846 net827 total_design.core.regFile.register\[1\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__a22o_1
XANTENNA__07111__B1 _02092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11994__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09237_ net336 _02565_ _04238_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__a21o_1
X_06449_ total_design.core.ctrl.instruction\[12\] net888 vssd1 vssd1 vccd1 vccd1 _02024_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_118_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09548__X _04780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09168_ _04364_ _04415_ net460 vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08119_ total_design.core.regFile.register\[30\]\[31\] net839 net803 total_design.core.regFile.register\[8\]\[31\]
+ _03610_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__a221o_1
X_09099_ _02286_ net319 vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__nand2_1
XANTENNA__10634__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11130_ _05386_ _05388_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__nand2_1
XANTENNA__07068__X _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold970 total_design.core.regFile.register\[3\]\[18\] vssd1 vssd1 vccd1 vccd1 net2286
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold981 total_design.core.regFile.register\[3\]\[29\] vssd1 vssd1 vccd1 vccd1 net2297
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ _05312_ _05315_ _05319_ _05313_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__or4b_1
Xhold992 total_design.core.regFile.register\[1\]\[20\] vssd1 vssd1 vccd1 vccd1 net2308
+ sky130_fd_sc_hd__dlygate4sd3_1
X_10012_ net184 net2758 net416 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__mux2_1
XANTENNA__07717__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11465__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12474__A1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11963_ net474 _05808_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__or2_4
XFILLER_0_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_83_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08142__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13702_ clknet_leaf_36_clk total_design.core.data_mem.stored_read_data\[9\] net1071
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10914_ _05145_ _05148_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__nand2_1
X_11894_ total_design.bus_full _01913_ _05772_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07350__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13633_ clknet_leaf_60_clk total_design.core.data_mem.data_write_adr_i\[5\] net1130
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[5\] sky130_fd_sc_hd__dfrtp_1
X_10845_ _05102_ _05103_ _05100_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__a21o_2
XFILLER_0_41_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13564_ clknet_leaf_41_clk total_design.core.data_mem.data_bus_i\[0\] net1092 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[0\] sky130_fd_sc_hd__dfrtp_1
X_10776_ total_design.core.data_bus_o\[22\] net695 vssd1 vssd1 vccd1 vccd1 _05035_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12515_ net976 total_design.core.instr_mem.instruction_i\[21\] vssd1 vssd1 vccd1
+ vccd1 _01712_ sky130_fd_sc_hd__and2b_1
X_13495_ clknet_leaf_161_clk _00962_ net1165 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08850__B1 _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12446_ net2559 net225 net346 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11737__B1 _05077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12377_ total_design.core.math.pc_val\[25\] net523 _01637_ _01638_ vssd1 vssd1 vccd1
+ vccd1 _01495_ sky130_fd_sc_hd__a22o_1
XANTENNA__10544__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07956__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11328_ net294 _05559_ _05544_ _05551_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__and4bb_1
X_14116_ clknet_leaf_100_clk _01296_ net1230 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output83_A net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11259_ _05419_ _05515_ _05508_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_157_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14047_ clknet_leaf_97_clk _01227_ net1245 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07169__B1 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07708__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06916__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_167_Right_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_74_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_35_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09330__A1 _02796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08133__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08470_ _01759_ _03800_ _03801_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_159_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07421_ total_design.core.ctrl.instruction\[16\] _02846_ total_design.core.ctrl.instruction\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wire308_X net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10719__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10228__B1 total_design.core.instr_fetch vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07352_ total_design.core.regFile.register\[4\]\[15\] net814 net769 total_design.core.regFile.register\[7\]\[15\]
+ net693 vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__a221o_1
X_06303_ _01854_ _01881_ _01866_ _01861_ _01858_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_169_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07283_ total_design.core.regFile.register\[22\]\[14\] net677 net631 total_design.core.regFile.register\[5\]\[14\]
+ _02802_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__a221o_1
XANTENNA__08841__B1 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09022_ _04268_ _04274_ net328 vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__mux2_1
X_06234_ total_design.core.data_adr_o\[19\] _01812_ net962 vssd1 vssd1 vccd1 vccd1
+ _01813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10962__B _05220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11728__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold200 total_design.lcd_display.row_1\[17\] vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold211 total_design.lcd_display.row_1\[71\] vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10454__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06165_ total_design.core.ctrl.instruction\[31\] vssd1 vssd1 vccd1 vccd1 _01748_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_14_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold222 total_design.lcd_display.row_1\[16\] vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold233 total_design.lcd_display.row_1\[77\] vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 total_design.core.math.pc_val\[0\] vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07947__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold255 total_design.lcd_display.row_1\[13\] vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold266 total_design.lcd_display.row_2\[76\] vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold277 total_design.lcd_display.row_1\[99\] vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold288 total_design.lcd_display.row_1\[44\] vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 total_design.lcd_display.row_1\[75\] vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout702 net703 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_2
X_09924_ net272 net2028 net424 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout713 _03917_ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1111_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout724 net725 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__buf_1
XANTENNA__12153__B1 _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout735 _02036_ vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_165_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout746 net748 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__clkbuf_2
Xfanout757 _02026_ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__buf_2
X_09855_ net258 net2389 net432 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__mux2_1
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout571_A _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06907__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 net770 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06887__B _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout779 net782 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_8
X_08806_ total_design.core.data_mem.data_cpu_i\[4\] _02335_ _02367_ _02388_ vssd1
+ vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__o2bb2a_1
X_09786_ net258 net2038 net440 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__mux2_1
X_06998_ total_design.core.regFile.register\[4\]\[9\] net622 net564 total_design.core.regFile.register\[3\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__a22o_1
XANTENNA__07580__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08737_ _02796_ _02845_ _02893_ _03992_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_65_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout836_A net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08124__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08668_ total_design.lcd_display.cnt_500hz\[13\] _03946_ net711 vssd1 vssd1 vccd1
+ vccd1 _03947_ sky130_fd_sc_hd__a21boi_1
XANTENNA__07332__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07619_ net551 net457 net288 vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__o21ai_2
XANTENNA__06686__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10629__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ total_design.data_in_BUS\[20\] net341 net715 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[20\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10219__A0 _04866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10630_ net282 net2485 net476 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06408__A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10561_ net246 net1869 net370 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ net899 _02993_ net522 vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13280_ clknet_leaf_193_clk _00747_ net1012 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10492_ net161 net2646 net378 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12231_ total_design.core.math.pc_val\[10\] total_design.core.program_count.imm_val_reg\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_20_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10364__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11687__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07399__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07938__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ _05767_ _05769_ _06012_ _06013_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__o211ai_2
XANTENNA__06143__A total_design.core.data_bus_o\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11113_ _05368_ _05369_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12093_ net126 net710 _05936_ _05950_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__o22a_1
X_11044_ _05302_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11990__Y _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_56_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11104__D1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12995_ clknet_leaf_8_clk _00462_ net1016 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08115__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11946_ _05745_ _05749_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07323__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06677__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10539__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11877_ _05757_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13616_ clknet_leaf_48_clk net1326 net1102 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10828_ _05072_ _05085_ _05061_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_138_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06429__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13547_ clknet_leaf_114_clk _01014_ net1202 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10759_ net961 _01773_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13478_ clknet_leaf_200_clk _00945_ net1002 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12429_ total_design.core.math.pc_val\[31\] net527 _01680_ _01684_ vssd1 vssd1 vccd1
+ vccd1 _01501_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10274__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09348__B _04588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07929__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07149__A _02666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07970_ total_design.core.regFile.register\[4\]\[28\] net814 net808 total_design.core.regFile.register\[5\]\[28\]
+ net692 vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06601__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12135__B1 _05826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06921_ total_design.core.regFile.register\[3\]\[7\] net866 net854 total_design.core.regFile.register\[16\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_143_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_0__f_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_09640_ net183 net2340 net455 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__mux2_1
X_06852_ total_design.core.regFile.register\[10\]\[6\] net617 net572 total_design.core.regFile.register\[17\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__a22o_1
XANTENNA__06500__B net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09571_ _04801_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__inv_2
X_06783_ total_design.core.ctrl.instruction\[25\] _02343_ vssd1 vssd1 vccd1 vccd1
+ _02344_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_47_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08522_ net2881 net342 _03872_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_136_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08453_ _03805_ _03806_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__nand2_1
XANTENNA__10449__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06668__A2 _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout152_A _05682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07404_ total_design.core.regFile.register\[16\]\[16\] net855 net761 total_design.core.regFile.register\[21\]\[16\]
+ _02930_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08384_ _03739_ _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07335_ total_design.core.regFile.register\[16\]\[15\] net635 _02861_ _02864_ vssd1
+ vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__a211o_1
XFILLER_0_116_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout417_A _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07266_ total_design.core.ctrl.instruction\[26\] net889 _02699_ _02799_ vssd1 vssd1
+ vccd1 vccd1 total_design.core.ctrl.imm_32\[14\] sky130_fd_sc_hd__a211o_1
XANTENNA__06515__X _02089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09005_ _04256_ _04257_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_115_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06217_ _01788_ _01791_ _01793_ _01795_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__or4b_1
XFILLER_0_115_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10184__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07197_ total_design.core.regFile.register\[15\]\[12\] net848 _02732_ _02733_ _02735_
+ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08162__B _02395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12374__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09973__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06148_ net1 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout786_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07250__C1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout510 net511 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12126__B1 _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout521 _01885_ vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_4
X_09907_ net194 net2538 net426 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__mux2_1
Xfanout543 net544 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout953_A _01911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout554 net555 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_2
XANTENNA_fanout574_X net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 _02094_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09542__B2 _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout576 _02089_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_4
X_09838_ net199 net2582 net436 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__mux2_1
Xfanout587 net588 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__buf_4
Xfanout598 net600 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07553__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06410__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09769_ net201 net2651 net444 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_38_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11800_ _03910_ _05702_ net713 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__o21bai_1
X_12780_ clknet_leaf_168_clk _00247_ net1158 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07305__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07522__A total_design.core.ctrl.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11731_ net1707 net957 net290 total_design.core.data_bus_o\[3\] vssd1 vssd1 vccd1
+ vccd1 _01359_ sky130_fd_sc_hd__a22o_1
XANTENNA__06659__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14450_ clknet_leaf_67_clk net1360 net1112 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11662_ _05665_ net1765 net131 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13401_ clknet_leaf_187_clk _00868_ net1028 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10613_ net207 net2377 net365 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11593_ _05677_ net1698 net137 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14381_ clknet_leaf_184_clk _01522_ net1039 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08805__B1 total_design.core.data_mem.data_cpu_i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13332_ clknet_leaf_142_clk _00799_ net1176 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10544_ net215 net2574 net373 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__mux2_1
XANTENNA__07084__A2 _01932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10094__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13263_ clknet_leaf_162_clk _00730_ net1153 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10475_ net232 net2279 net380 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11168__A1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12214_ total_design.core.math.pc_val\[8\] total_design.core.program_count.imm_val_reg\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__or2_1
XANTENNA__11985__Y _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13194_ clknet_leaf_24_clk _00661_ net1108 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12145_ total_design.lcd_display.row_2\[39\] _05847_ _05850_ total_design.lcd_display.row_2\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12117__B1 _05832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12076_ total_design.lcd_display.row_1\[52\] _05840_ _05849_ total_design.lcd_display.row_2\[52\]
+ _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__a221o_1
XANTENNA__08336__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11027_ net351 _05281_ _05285_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__a21o_1
XANTENNA__09533__A1 _03234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06898__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11653__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12978_ clknet_leaf_146_clk _00445_ net1177 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11929_ total_design.keypad0.key_out\[9\] net529 net475 total_design.keypad0.key_out\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10269__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08247__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09049__A0 _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10793__A total_design.core.data_bus_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07120_ _02655_ _02657_ _02659_ _02661_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__or4_1
XFILLER_0_70_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07075__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07051_ total_design.core.regFile.register\[15\]\[10\] net604 net569 total_design.core.regFile.register\[17\]\[10\]
+ _02595_ vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a221o_1
XANTENNA__11401__B _05652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06822__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09793__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XANTENNA__09221__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_162_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07953_ total_design.core.regFile.register\[7\]\[27\] net653 net605 total_design.core.regFile.register\[15\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06904_ total_design.core.regFile.register\[23\]\[7\] net681 net616 total_design.core.regFile.register\[10\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__a22o_1
X_07884_ total_design.core.regFile.register\[8\]\[26\] net803 _03382_ _03383_ _03385_
+ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07535__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ net465 _04811_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__nor2_1
X_06835_ _02391_ _02392_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__or2_1
XANTENNA__11416__X _05675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__S net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09554_ _04784_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__inv_2
X_06766_ total_design.core.regFile.register\[16\]\[4\] net632 net581 total_design.core.regFile.register\[6\]\[4\]
+ _02327_ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__a221o_1
XFILLER_0_167_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09033__S net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08505_ _03855_ _03856_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10179__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06697_ _02263_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[3\]
+ sky130_fd_sc_hd__inv_2
X_09485_ _04714_ _04719_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__or2_4
XANTENNA__06229__Y _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout155_X net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout534_A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08157__B _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09968__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08436_ _03760_ _03789_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08367_ total_design.keypad0.key_out\[1\] total_design.keypad0.key_out\[4\] vssd1
+ vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout701_A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout322_X net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07318_ total_design.core.ctrl.instruction\[27\] net887 _02699_ _02848_ vssd1 vssd1
+ vccd1 vccd1 total_design.core.ctrl.imm_32\[15\] sky130_fd_sc_hd__a211o_1
X_08298_ net1455 net941 _03683_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[6\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12407__B _03559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08604__C net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07249_ total_design.core.regFile.register\[15\]\[13\] net846 net759 total_design.core.regFile.register\[21\]\[13\]
+ _02784_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06813__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1231_X net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10260_ net166 net2253 net503 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ net269 net1945 net389 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__mux2_1
XANTENNA__10642__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07517__A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout340 net341 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_2
Xfanout351 _05043_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_2
Xfanout362 net363 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_8
X_13950_ clknet_leaf_97_clk _01130_ net1244 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[32\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout373 _05012_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_8
Xfanout384 _05009_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout395 net396 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_8
X_12901_ clknet_leaf_116_clk _00368_ net1203 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13881_ clknet_leaf_38_clk total_design.core.ctrl.imm_32\[20\] net1080 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11473__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09451__B _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12832_ clknet_leaf_194_clk _00299_ net1011 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12763_ clknet_leaf_149_clk _00230_ net1174 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10089__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09878__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14502_ clknet_leaf_33_clk _01569_ net1070 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[30\]
+ sky130_fd_sc_hd__dfrtp_4
X_11714_ net19 net934 net877 net2184 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__o22a_1
XFILLER_0_167_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12694_ clknet_leaf_155_clk _00161_ net1138 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14433_ clknet_leaf_34_clk total_design.core.data_out_INSTR\[28\] net1069 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[28\] sky130_fd_sc_hd__dfrtp_1
X_11645_ _05643_ net1846 net133 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07057__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14364_ clknet_leaf_154_clk _01505_ net1136 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_11576_ _05612_ net1671 net141 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__mux2_1
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
Xinput37 gpio_in[32] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
XFILLER_0_25_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13315_ clknet_leaf_16_clk _00782_ net1024 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06804__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10527_ net286 net1877 net374 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__mux2_1
X_14295_ clknet_leaf_95_clk _01471_ net1256 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.lcd_rs
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13246_ clknet_leaf_167_clk _00713_ net1155 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10458_ net167 net1927 net383 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08811__A _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11648__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10552__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13177_ clknet_leaf_195_clk _00644_ net1010 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10389_ net176 net1917 net487 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__mux2_1
X_12128_ total_design.lcd_display.row_1\[94\] _05812_ _05826_ total_design.lcd_display.row_1\[22\]
+ _05983_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__a221o_1
XFILLER_0_165_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08309__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12059_ total_design.lcd_display.row_1\[75\] _05816_ _05909_ _05916_ _05917_ vssd1
+ vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_88_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10788__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06620_ total_design.core.regFile.register\[29\]\[2\] net926 net947 net910 vssd1
+ vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__and4_1
XFILLER_0_88_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13501__RESET_B net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06551_ total_design.core.regFile.register\[10\]\[1\] net920 net916 net913 vssd1
+ vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__and4_1
XFILLER_0_158_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09788__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09270_ net316 _04302_ _04513_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_103_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06482_ net745 net730 net724 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__and3_4
XANTENNA__07296__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09690__B1 _03559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08221_ net1368 net545 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[4\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_7_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08152_ net553 total_design.core.data_mem.data_cpu_i\[31\] total_design.core.ctrl.imm_32\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__a21oi_4
XANTENNA__12041__A2 _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09442__B1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07103_ _02644_ _02645_ _02643_ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_151_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08083_ total_design.core.regFile.register\[0\]\[30\] net876 _03562_ _03576_ vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[30\] sky130_fd_sc_hd__o22a_4
XFILLER_0_141_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_9_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07034_ total_design.core.regFile.register\[5\]\[9\] net808 _02580_ _02581_ vssd1
+ vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__a211o_1
XANTENNA__11558__S net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10462__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11552__A1 _05630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07756__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1024_A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07220__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08985_ net336 _02515_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout484_A _05007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06598__D net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ total_design.core.regFile.register\[3\]\[27\] net867 net843 total_design.core.regFile.register\[25\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__a22o_1
XANTENNA__07508__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07867_ net553 total_design.core.data_mem.data_cpu_i\[25\] total_design.core.ctrl.imm_32\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout651_A _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout749_A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09606_ _04670_ _04687_ _04832_ _04834_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06818_ total_design.core.regFile.register\[3\]\[5\] net868 net856 total_design.core.regFile.register\[16\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_27_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08168__A _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07798_ net553 net307 _03179_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11068__B1 _05184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09537_ net465 _04174_ _04177_ _04767_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a31o_1
X_06749_ _01739_ net949 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1181_X net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout537_X net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09130__C1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09468_ _03088_ _04701_ _04702_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07287__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08419_ total_design.keypad0.key_out\[6\] _03715_ vssd1 vssd1 vccd1 vccd1 _03774_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10637__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09399_ _02868_ _02889_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11430_ net1515 _05667_ net157 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12032__A2 _05814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11361_ net303 _05475_ _05614_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07995__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13100_ clknet_leaf_165_clk _00567_ net1165 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10312_ net221 net2433 net494 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11292_ net248 _05549_ _05543_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__o21ba_1
X_14080_ clknet_leaf_110_clk _01260_ net1227 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11468__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09197__C1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10243_ net231 net2048 net503 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__mux2_1
X_13031_ clknet_leaf_19_clk _00498_ net1049 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10372__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__A1 _05612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1102 net1104 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_4
X_10174_ net209 net2234 net395 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__mux2_1
Xfanout1113 net1116 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__clkbuf_4
Xfanout1124 net1134 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__clkbuf_4
Xfanout1135 net39 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__buf_4
Xfanout1146 net1149 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12099__A2 _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1157 net1163 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__clkbuf_4
Xfanout170 _04929_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1168 net1172 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__clkbuf_2
Xfanout181 net184 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_2
Xfanout1179 net1181 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__clkbuf_4
Xfanout192 _04822_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_2
X_13933_ clknet_leaf_92_clk _01113_ net1262 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13864_ clknet_leaf_65_clk total_design.core.ctrl.imm_32\[3\] net1124 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06722__A1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12815_ clknet_leaf_146_clk _00282_ net1178 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13795_ clknet_leaf_76_clk total_design.core.data_mem.data_cpu_i\[4\] net1213 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10806__B1 _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12746_ clknet_leaf_23_clk _00213_ net1055 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10547__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12677_ clknet_leaf_118_clk _00144_ net1160 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10774__C _05028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14416_ clknet_leaf_36_clk total_design.core.data_out_INSTR\[11\] net1071 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11628_ _05663_ net1757 net134 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06326__A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12023__A2 _05812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14347_ clknet_leaf_44_clk _00034_ net1087 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11559_ _05626_ net1662 net143 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__mux2_1
Xhold607 total_design.core.regFile.register\[5\]\[6\] vssd1 vssd1 vccd1 vccd1 net1923
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold618 total_design.core.regFile.register\[7\]\[17\] vssd1 vssd1 vccd1 vccd1 net1934
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09196__X _04443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold629 total_design.core.regFile.register\[16\]\[3\] vssd1 vssd1 vccd1 vccd1 net1945
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14278_ net987 _01454_ net1082 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[7\]
+ sky130_fd_sc_hd__dfrtp_4
Xmax_cap348 _05835_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_4
XANTENNA__07450__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10282__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13229_ clknet_leaf_5_clk _00696_ net1022 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06332__Y _01911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11534__A1 _05679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08260__B net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1092 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07738__B1 _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07157__A total_design.core.ctrl.instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_97_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1307 total_design.core.regFile.register\[6\]\[13\] vssd1 vssd1 vccd1 vccd1 net2623
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1318 total_design.data_in_BUS\[31\] vssd1 vssd1 vccd1 vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
X_08770_ total_design.core.data_mem.data_cpu_i\[31\] net305 vssd1 vssd1 vccd1 vccd1
+ _04025_ sky130_fd_sc_hd__or2_1
Xhold1329 total_design.core.regFile.register\[25\]\[20\] vssd1 vssd1 vccd1 vccd1 net2645
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07444__X _02968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07721_ _03229_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__inv_2
X_07652_ total_design.core.regFile.register\[30\]\[21\] net660 net602 total_design.core.regFile.register\[31\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07910__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06603_ total_design.core.regFile.register\[12\]\[1\] _02092_ _02160_ _02163_ _02168_
+ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_157_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07583_ total_design.core.regFile.register\[23\]\[20\] net678 net593 total_design.core.regFile.register\[8\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_122_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09322_ net506 _04563_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__and2_1
X_06534_ net906 net888 _02028_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_122_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07269__A2 _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11065__A3 _05064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09253_ _02565_ _02584_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06465_ _01924_ net901 _02018_ total_design.core.ctrl.instruction\[16\] _01741_ vssd1
+ vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__o311a_1
XANTENNA__10457__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08204_ total_design.core.data_mem.data_read_adr_reg\[25\] total_design.core.data_mem.data_read_adr_reg\[24\]
+ total_design.core.data_mem.data_read_adr_reg\[27\] total_design.core.data_mem.data_read_adr_reg\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__or4_1
X_09184_ _02492_ net703 _04430_ net534 vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__a211o_1
XANTENNA__12014__A2 _05829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06396_ net923 _01950_ net908 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_170_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06229__B1 net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08135_ total_design.core.regFile.register\[29\]\[31\] net656 net617 total_design.core.regFile.register\[10\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1141_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14529__1301 vssd1 vssd1 vccd1 vccd1 net1301 _14529__1301/LO sky130_fd_sc_hd__conb_1
XANTENNA__07977__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1239_A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ total_design.core.regFile.register\[3\]\[30\] net868 net785 total_design.core.regFile.register\[2\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__a22o_1
XANTENNA__07441__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07017_ _02564_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10192__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09266__B net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08170__B _02796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07729__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1027_X net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09981__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout866_A _01941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_X net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ net473 _02770_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__or2_1
X_07919_ _03323_ _03327_ _03372_ _03418_ _03371_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__a311oi_1
XANTENNA_fanout654_X net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08899_ net337 _02182_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__nor2_1
X_10930_ _05156_ _05159_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__nor2_1
XANTENNA__07901__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861_ _05118_ _05119_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout821_X net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout919_X net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ clknet_leaf_136_clk _00067_ net1179 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13580_ clknet_leaf_27_clk total_design.core.data_mem.data_bus_i\[16\] net1073 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[16\] sky130_fd_sc_hd__dfrtp_1
X_10792_ total_design.core.data_bus_o\[10\] total_design.core.data_bus_o\[6\] total_design.core.data_bus_o\[5\]
+ total_design.core.data_bus_o\[4\] vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__and4b_1
XFILLER_0_66_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12531_ net977 total_design.core.instr_mem.instruction_i\[29\] vssd1 vssd1 vccd1
+ vccd1 _01720_ sky130_fd_sc_hd__and2b_1
XANTENNA__10367__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12005__A2 _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12462_ net2742 net162 net345 vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__mux2_1
XANTENNA__07680__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14201_ clknet_leaf_80_clk _01381_ net1222 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
X_11413_ _05670_ _05671_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12393_ net991 _04886_ net894 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11764__A1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14132_ clknet_leaf_99_clk _01312_ net1229 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11344_ _05449_ _05453_ _05451_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__a21o_1
XANTENNA__07432__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14063_ clknet_leaf_97_clk _01243_ net1245 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[81\]
+ sky130_fd_sc_hd__dfrtp_1
X_11275_ _05532_ _05533_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__nand2_1
XANTENNA__11516__A1 _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09891__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13014_ clknet_leaf_156_clk _00481_ net1142 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10226_ _04966_ net391 _05000_ vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10157_ net276 net2509 net395 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__mux2_1
XANTENNA__09463__Y _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold4 total_design.core.data_mem.data_read_adr_reg\[2\] vssd1 vssd1 vccd1 vccd1 net1320
+ sky130_fd_sc_hd__dlygate4sd3_1
X_10088_ net245 net2447 net402 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08145__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13916_ clknet_leaf_99_clk _01096_ net1227 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07499__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12492__A2 total_design.core.ctrl.instruction\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13847_ clknet_leaf_48_clk _01055_ net1102 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11661__S net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13778_ clknet_leaf_48_clk total_design.core.data_mem.stored_data_adr\[21\] net1098
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[21\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13799__D total_design.core.data_mem.data_cpu_i\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_127_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12729_ clknet_leaf_196_clk _00196_ net1009 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10277__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08255__B net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06250_ _01771_ _01828_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06181_ total_design.core.mem_ctrl.state\[1\] total_design.core.mem_ctrl.state\[2\]
+ total_design.core.mem_ctrl.state\[0\] vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__or3b_4
XFILLER_0_81_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold404 net71 vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11755__B2 total_design.core.data_bus_o\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold415 total_design.core.math.pc_val\[12\] vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold426 net68 vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold437 net100 vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold448 total_design.core.math.pc_val\[1\] vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 total_design.lcd_display.row_2\[34\] vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09940_ net199 net1952 net423 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__mux2_1
XANTENNA__06631__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11507__A1 _05652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06503__B net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout906 _02014_ vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09871_ net201 net2703 net431 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__mux2_1
Xfanout917 _01935_ vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__buf_2
Xfanout928 _01925_ vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__buf_2
Xfanout939 _03675_ vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_74_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _04061_ _04076_ _04068_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_146_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09814__B total_design.core.ctrl.instruction\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 total_design.core.regFile.register\[6\]\[14\] vssd1 vssd1 vccd1 vccd1 net2420
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 total_design.core.regFile.register\[7\]\[5\] vssd1 vssd1 vccd1 vccd1 net2431
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 total_design.core.regFile.register\[15\]\[26\] vssd1 vssd1 vccd1 vccd1 net2442
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 total_design.core.regFile.register\[14\]\[16\] vssd1 vssd1 vccd1 vccd1 net2453
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11408__Y _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08753_ _04006_ _04007_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1148 total_design.core.regFile.register\[8\]\[16\] vssd1 vssd1 vccd1 vccd1 net2464
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout182_A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08136__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1159 total_design.core.regFile.register\[16\]\[0\] vssd1 vssd1 vccd1 vccd1 net2475
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_124_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07704_ total_design.core.regFile.register\[15\]\[22\] net605 net583 total_design.core.regFile.register\[6\]\[22\]
+ _03212_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08684_ net1406 _03960_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07635_ total_design.core.regFile.register\[1\]\[21\] net828 net820 total_design.core.regFile.register\[17\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11571__S net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout447_A _04189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12235__A2 _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07566_ total_design.core.data_mem.data_cpu_i\[19\] vssd1 vssd1 vccd1 vccd1 _03083_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_137_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06518__X _02092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09305_ _02746_ net702 vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__nand2_1
X_06517_ net745 net736 net728 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__and3_4
XFILLER_0_152_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07497_ total_design.core.regFile.register\[9\]\[18\] net850 net802 total_design.core.regFile.register\[8\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout614_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09976__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09236_ _02589_ net702 _04480_ net534 vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__a211o_1
X_06448_ _01735_ _01919_ _02012_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__and3_1
XANTENNA__07662__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06870__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06379_ total_design.core.regFile.register\[25\]\[0\] net927 net913 net910 vssd1
+ vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09167_ _04143_ _04147_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1144_X net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11746__B2 total_design.core.data_bus_o\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08118_ total_design.core.regFile.register\[3\]\[31\] net867 net795 total_design.core.regFile.register\[11\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_3_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ net269 net2322 net453 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout983_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ total_design.core.regFile.register\[15\]\[29\] net604 net581 total_design.core.regFile.register\[6\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold960 total_design.core.regFile.register\[31\]\[19\] vssd1 vssd1 vccd1 vccd1 net2276
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06413__B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold971 total_design.core.regFile.register\[3\]\[17\] vssd1 vssd1 vccd1 vccd1 net2287
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ _05317_ _05318_ _05316_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__a21oi_1
Xhold982 total_design.core.regFile.register\[27\]\[29\] vssd1 vssd1 vccd1 vccd1 net2298
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold993 total_design.core.regFile.register\[9\]\[5\] vssd1 vssd1 vccd1 vccd1 net2309
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ net188 net2659 net416 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout869_X net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10650__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06700__Y _02266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08127__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11962_ _05733_ _05823_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__and2_1
XANTENNA__11682__A0 _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13701_ clknet_leaf_38_clk total_design.core.data_mem.stored_read_data\[8\] net1079
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10913_ _05145_ _05170_ _05146_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__a21bo_1
XANTENNA__06689__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11893_ wishbone.curr_state\[0\] _01912_ _01910_ vssd1 vssd1 vccd1 vccd1 _05772_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11481__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13632_ clknet_leaf_60_clk total_design.core.data_mem.data_write_adr_i\[4\] net1130
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10844_ _05092_ _05096_ _05098_ _05088_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13563_ clknet_leaf_146_clk _01030_ net1177 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10097__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10775_ total_design.core.data_bus_o\[25\] net700 vssd1 vssd1 vccd1 vccd1 _05034_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09886__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12514_ net976 total_design.core.ctrl.instruction\[20\] net882 _01711_ vssd1 vssd1
+ vccd1 vccd1 _01559_ sky130_fd_sc_hd__a22o_1
XANTENNA__11988__Y _05850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07653__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13494_ clknet_leaf_155_clk _00961_ net1137 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08850__A1 total_design.core.ctrl.instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12445_ net2844 net232 net347 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07405__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12376_ net900 _03375_ net523 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__a21oi_1
X_14115_ clknet_leaf_89_clk _01295_ net1261 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06613__B1 total_design.core.ctrl.imm_32\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11327_ _05582_ _05585_ net294 vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07419__B _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ clknet_leaf_100_clk _01226_ net1229 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_11258_ _05427_ _05429_ _05516_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11656__S net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10209_ _04680_ net2672 net389 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10560__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11189_ _05442_ _05447_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08118__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11673__A0 _05636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14528__1300 vssd1 vssd1 vccd1 vccd1 net1300 _14528__1300/LO sky130_fd_sc_hd__conb_1
XFILLER_0_159_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10796__A _01885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07420_ total_design.core.ctrl.instruction\[16\] total_design.core.ctrl.instruction\[17\]
+ _02846_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__or3_1
XANTENNA__07892__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10228__A1 total_design.core.ctrl.instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07351_ total_design.core.regFile.register\[21\]\[15\] net761 _02879_ _02880_ vssd1
+ vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10779__A2 total_design.core.data_bus_o\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06302_ _01875_ _01879_ _01808_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09796__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07282_ total_design.core.regFile.register\[29\]\[14\] net658 net566 total_design.core.regFile.register\[12\]\[14\]
+ _02804_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06233_ total_design.core.instr_mem.instruction_adr_i\[19\] total_design.core.instr_mem.instruction_adr_stored\[19\]
+ net981 vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__mux2_1
XANTENNA__06217__C _01793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09021_ _04270_ _04273_ net467 vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06852__B1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11728__A1 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06164_ net967 vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__inv_2
Xhold201 total_design.lcd_display.row_1\[10\] vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 total_design.lcd_display.row_1\[116\] vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 total_design.lcd_display.row_1\[85\] vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold234 total_design.lcd_display.row_1\[70\] vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold245 total_design.lcd_display.row_1\[121\] vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold256 total_design.lcd_display.row_1\[41\] vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 total_design.lcd_display.row_1\[102\] vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 total_design.lcd_display.row_1\[114\] vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09923_ net260 net2380 net424 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold289 total_design.lcd_display.row_1\[48\] vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout703 _04204_ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__buf_2
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout714 net716 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11566__S net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 _02048_ vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout736 net737 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__buf_2
X_09854_ net280 net2087 net430 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__mux2_1
XANTENNA__10470__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout747 net748 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__clkbuf_2
Xfanout758 _02004_ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1104_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout769 net770 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_4
X_08805_ _02263_ _02286_ total_design.core.data_mem.data_cpu_i\[4\] _02335_ vssd1
+ vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__o2bb2a_1
X_09785_ net281 net2700 net438 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout564_A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06997_ total_design.core.regFile.register\[23\]\[9\] net680 net572 total_design.core.regFile.register\[17\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__a22o_1
XANTENNA__09306__C1 _04105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_192_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ _02640_ _02695_ _02746_ _03991_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__and4_1
XANTENNA__11664__A0 _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09321__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08667_ _03946_ net711 _03945_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout829_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07618_ net457 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[20\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__07883__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08598_ total_design.data_in_BUS\[19\] net341 net715 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[19\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_166_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08607__C net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ total_design.core.regFile.register\[16\]\[19\] net855 net832 total_design.core.regFile.register\[31\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06408__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_X net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07635__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10560_ net284 net2564 net370 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_130_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06843__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ net316 _04183_ _04191_ _04464_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__o211a_1
XANTENNA__10645__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10491_ net166 net2427 net379 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12230_ net902 _02640_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12161_ _06012_ _06013_ _05767_ _05769_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_145_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11112_ _05366_ _05367_ _05370_ _05368_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_9_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09735__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12092_ _05945_ _05949_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__or2_1
Xhold790 total_design.core.regFile.register\[18\]\[30\] vssd1 vssd1 vccd1 vccd1 net2106
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11476__S net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ _05236_ _05238_ _05301_ _05056_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_120_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10380__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10155__A0 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06359__C1 total_design.core.ctrl.instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07020__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11104__C1 _05064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ clknet_leaf_126_clk _00461_ net1193 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11655__A0 _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1490 total_design.core.regFile.register\[24\]\[14\] vssd1 vssd1 vccd1 vccd1 net2806
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11945_ _05732_ _05742_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__nand2_4
XFILLER_0_8_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07261__Y _02796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11876_ net995 net902 vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__nor2_2
XANTENNA__07874__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13615_ clknet_leaf_49_clk net1343 net1103 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10827_ _05076_ _05085_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12080__B1 _05848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13546_ clknet_leaf_25_clk _01013_ net1106 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10758_ net1861 _05019_ _01775_ vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08814__A total_design.core.data_mem.data_cpu_i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_125_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10555__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13477_ clknet_leaf_117_clk _00944_ net1212 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10689_ net165 net2126 net363 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11882__A2_N _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12428_ net902 _03646_ _05760_ _01683_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__a22oi_1
XANTENNA__06334__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12359_ total_design.core.math.pc_val\[24\] net988 vssd1 vssd1 vccd1 vccd1 _01622_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07717__X _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14029_ clknet_leaf_92_clk _01209_ net1258 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10290__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06920_ total_design.core.regFile.register\[31\]\[7\] net831 net822 total_design.core.regFile.register\[17\]\[7\]
+ _02473_ vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_71_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11894__A0 total_design.bus_full vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ total_design.core.regFile.register\[21\]\[6\] net599 net579 total_design.core.regFile.register\[27\]\[6\]
+ _02407_ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_160_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09570_ _04799_ _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_160_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06782_ _02149_ _02312_ _02028_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__a21o_1
X_08521_ _03856_ _03858_ _03870_ _03871_ _03767_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__a311o_1
XANTENNA__11646__A0 _05645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11415__A _05609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ _03799_ _03804_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07403_ total_design.core.regFile.register\[31\]\[16\] net833 net812 total_design.core.regFile.register\[23\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__a22o_1
X_08383_ total_design.keypad0.key_out\[8\] _03726_ _03727_ vssd1 vssd1 vccd1 vccd1
+ _03740_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_9_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout145_A net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07078__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12071__B1 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07334_ total_design.core.regFile.register\[22\]\[15\] net676 _02862_ _02863_ vssd1
+ vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__a211o_1
XANTENNA__07617__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10465__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07265_ _02797_ _02798_ net722 vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08290__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1054_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09004_ net471 net308 vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06216_ total_design.core.data_adr_o\[25\] _01794_ net961 vssd1 vssd1 vccd1 vccd1
+ _01795_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_115_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07196_ total_design.core.regFile.register\[11\]\[12\] net794 _02720_ _02734_ vssd1
+ vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__a211o_1
XFILLER_0_103_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06147_ total_design.key_confirm vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1221_A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08042__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07250__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout500 net503 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_6
Xfanout511 net512 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout779_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout522 net525 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__buf_2
X_09906_ net200 net2512 net428 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__mux2_1
Xfanout533 net536 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_4
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07538__D1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout555 _02107_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_2
Xfanout566 _02092_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07002__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ net203 net2319 net436 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__mux2_1
Xfanout577 net580 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_8
Xfanout588 _02083_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout567_X net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout599 net600 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__buf_4
XANTENNA_fanout946_A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06410__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09768_ net205 net2749 net442 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08719_ _03950_ _03975_ _03979_ vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__nor3_1
X_09699_ _04922_ _04923_ net450 vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_68_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11730_ net95 net960 net293 net2223 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07856__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11661_ _05663_ net1804 net132 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__mux2_1
XANTENNA__09058__A1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ clknet_leaf_133_clk _00867_ net1195 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ net209 net2547 net366 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07069__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12062__B1 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07608__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14380_ clknet_leaf_161_clk _01521_ net1151 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11592_ _05626_ net1685 net139 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13331_ clknet_leaf_181_clk _00798_ net1042 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06816__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10375__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10543_ net221 net2373 net375 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12156__A _05823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13262_ clknet_leaf_189_clk _00729_ net1030 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10474_ net230 net2265 net380 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__mux2_1
XANTENNA__06154__A total_design.core.ctrl.instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11168__A2 _05184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12213_ total_design.core.math.pc_val\[8\] total_design.core.program_count.imm_val_reg\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08033__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ clknet_leaf_177_clk _00660_ net1046 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_92_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12144_ _05991_ _05993_ _05996_ _05998_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__or4_1
XANTENNA__07241__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06441__X _02016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12075_ total_design.lcd_display.row_1\[4\] _05830_ _05841_ total_design.lcd_display.row_1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11026_ _05056_ _05283_ _05284_ _05282_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__a31o_2
XANTENNA__09533__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_2__f_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08809__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11628__A0 _05663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12977_ clknet_leaf_148_clk _00444_ net1146 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11928_ total_design.keypad0.key_out\[8\] net530 net475 total_design.keypad0.key_out\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__a22o_1
XANTENNA__10300__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06329__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11859_ _05737_ _05743_ total_design.lcd_display.currentState\[5\] vssd1 vssd1 vccd1
+ vccd1 _05744_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08792__A_N total_design.core.data_mem.data_cpu_i\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06807__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13529_ clknet_leaf_196_clk _00996_ net1009 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10285__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08263__B net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07050_ total_design.core.regFile.register\[2\]\[10\] net636 net620 total_design.core.regFile.register\[4\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a22o_1
XANTENNA__07480__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11401__C _05655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XANTENNA__08024__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07232__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09375__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07952_ total_design.core.regFile.register\[14\]\[27\] net625 net586 total_design.core.regFile.register\[28\]\[27\]
+ _03450_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09662__X _04889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06903_ total_design.core.regFile.register\[29\]\[7\] net655 net589 total_design.core.regFile.register\[1\]\[7\]
+ _02456_ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a221o_1
X_07883_ total_design.core.regFile.register\[10\]\[26\] net836 net777 total_design.core.regFile.register\[22\]\[26\]
+ _03384_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__a221o_1
X_09622_ net332 _04769_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__nor2_1
X_06834_ _02392_ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__inv_2
X_09553_ _03207_ _03226_ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_108_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06765_ total_design.core.regFile.register\[5\]\[4\] net628 net604 total_design.core.regFile.register\[15\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout262_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08504_ _03834_ _03854_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07299__B1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09484_ total_design.core.ctrl.instruction\[19\] net887 net754 total_design.core.data_cpu_o\[19\]
+ _04718_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__a221o_1
XANTENNA__07838__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06696_ total_design.core.regFile.register\[0\]\[3\] net875 _02248_ _02262_ vssd1
+ vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_77_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08435_ _03760_ _03789_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout148_X net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1171_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12044__B1 _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08366_ total_design.data_in_BUS\[2\] net512 _01904_ vssd1 vssd1 vccd1 vccd1 _03724_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07317_ _02846_ _02847_ net721 vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__a21oi_1
X_08297_ total_design.core.data_mem.data_write_adr_reg\[6\] net549 net541 total_design.core.data_mem.data_read_adr_reg\[6\]
+ net945 vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__a221o_1
XANTENNA__08173__B _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13__f_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07248_ total_design.core.regFile.register\[28\]\[13\] net853 net783 total_design.core.regFile.register\[2\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout896_A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07179_ total_design.core.regFile.register\[0\]\[12\] net682 _02714_ _02717_ vssd1
+ vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__o22a_4
XANTENNA__07223__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ net276 net1990 net389 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06421__B net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout330 net331 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_2
Xfanout341 net343 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_2
Xfanout352 _05043_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_2
XANTENNA__09515__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout851_X net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout363 net364 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_8
Xfanout374 _05012_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_4
Xfanout385 net388 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_6
XANTENNA_fanout949_X net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_6
X_12900_ clknet_leaf_108_clk _00367_ net1223 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13880_ clknet_leaf_26_clk total_design.core.ctrl.imm_32\[19\] net1080 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[19\] sky130_fd_sc_hd__dfrtp_1
X_12831_ clknet_leaf_183_clk _00298_ net1039 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12762_ clknet_leaf_134_clk _00229_ net1196 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14501_ clknet_leaf_37_clk _01568_ net1076 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_51_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11713_ net18 net936 net879 net2477 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13800__RESET_B net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12693_ clknet_leaf_160_clk _00160_ net1142 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14432_ clknet_leaf_34_clk total_design.core.data_out_INSTR\[27\] net1069 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[27\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12035__B1 _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11644_ _05648_ net1712 net134 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06436__X total_design.core.data_mem.data_cpu_i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14363_ clknet_leaf_157_clk _01504_ net1044 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11575_ _05609_ net1715 net143 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__mux2_1
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_94_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput38 gpio_in[33] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09894__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13314_ clknet_leaf_127_clk _00781_ net1192 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09747__X _04969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07462__B1 _01992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10526_ _04982_ net532 vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__nand2_8
XFILLER_0_165_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14294_ clknet_leaf_91_clk _01470_ net1263 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13245_ clknet_leaf_10_clk _00712_ net1020 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10457_ net171 net2771 net381 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__mux2_1
XANTENNA__08006__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08811__B net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13176_ clknet_leaf_133_clk _00643_ net1195 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10388_ net181 net2508 net486 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__mux2_1
XANTENNA__06612__A _02182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ total_design.lcd_display.row_1\[6\] _05830_ _05841_ total_design.lcd_display.row_1\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__a22o_1
XANTENNA__09506__A2 _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12058_ total_design.lcd_display.row_1\[83\] _05815_ _05827_ total_design.lcd_display.row_1\[35\]
+ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__a22o_1
XANTENNA__11664__S net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ _05056_ _05267_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__nand2_1
XANTENNA__09642__B _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10788__B total_design.core.data_bus_o\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08258__B net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06740__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06550_ total_design.core.regFile.register\[25\]\[1\] net925 net913 net909 vssd1
+ vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__and4_1
XFILLER_0_88_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06481_ net746 net728 net723 vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__and3_1
XANTENNA__13541__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09690__B2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08220_ net1366 net545 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[3\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_172_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12026__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08151_ total_design.core.regFile.register\[0\]\[31\] net684 _03635_ _03641_ vssd1
+ vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_15_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09442__A1 total_design.core.data_cpu_o\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06506__B net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07102_ net896 _02019_ _02022_ _01748_ vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_151_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08082_ total_design.core.regFile.register\[21\]\[30\] net761 _03563_ _03564_ _03575_
+ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_114_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07033_ total_design.core.regFile.register\[9\]\[9\] net852 net796 total_design.core.regFile.register\[11\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07618__A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08984_ net469 _02468_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__nor2_1
XANTENNA__09392__X _04631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07935_ total_design.core.regFile.register\[31\]\[27\] net832 net768 total_design.core.regFile.register\[7\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__a22o_1
XANTENNA__11574__S net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07866_ total_design.core.regFile.register\[0\]\[25\] net684 _03362_ _03368_ vssd1
+ vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_127_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09605_ _03373_ net509 net448 _03372_ _04833_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06817_ total_design.core.regFile.register\[6\]\[5\] net765 _02376_ vssd1 vssd1 vccd1
+ vccd1 _02377_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07797_ net307 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[24\]
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout644_A _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06731__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09979__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ _04174_ _04177_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__nand2_1
X_06748_ _01930_ _02149_ _02020_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09467_ _03088_ _04701_ net706 vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06679_ total_design.core.regFile.register\[8\]\[3\] net803 net799 total_design.core.regFile.register\[29\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout811_A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout909_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12017__B1 _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08418_ _03771_ _03772_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__or2_1
XFILLER_0_163_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07692__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09398_ net225 net2848 net456 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__mux2_1
XANTENNA__07092__A_N _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ total_design.core.mem_ctrl.next_next_data_read _01774_ vssd1 vssd1 vccd1
+ vccd1 _03709_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06416__B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11360_ _05471_ _05606_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06798__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10311_ net225 net2370 net494 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__mux2_1
XANTENNA__10653__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291_ net248 _05549_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13030_ clknet_leaf_195_clk _00497_ net1008 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10242_ net236 net2652 net502 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__mux2_1
XANTENNA__09736__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1103 net1104 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__clkbuf_2
X_10173_ net216 net2598 net394 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1114 net1116 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__buf_2
Xfanout1125 net1128 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__clkbuf_4
Xfanout1136 net1144 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input38_A gpio_in[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1148 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__clkbuf_4
Xfanout160 _05676_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_2
Xfanout1158 net1163 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__buf_2
XANTENNA__11484__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_137_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout171 _04929_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1169 net1171 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06970__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout182 net184 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_2
X_13932_ clknet_leaf_98_clk _01112_ net1244 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[78\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout193 net196 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07263__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06183__A0 total_design.bus_full vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13863_ clknet_leaf_66_clk total_design.core.ctrl.imm_32\[2\] net1122 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06722__A2 _02263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11059__A1 total_design.core.data_bus_o\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12814_ clknet_leaf_187_clk _00281_ net1031 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09889__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13794_ clknet_leaf_76_clk total_design.core.data_mem.data_cpu_i\[3\] net1214 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10806__A1 total_design.core.data_bus_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ clknet_leaf_4_clk _00212_ net1023 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07683__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ clknet_leaf_128_clk _00143_ net1191 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_146_Left_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ clknet_leaf_38_clk total_design.core.data_out_INSTR\[10\] net1078 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[10\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _05627_ net1722 net136 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06326__B _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14346_ clknet_leaf_46_clk _00033_ net1086 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07435__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ _05624_ net1797 net144 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire561 _03670_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_1
XFILLER_0_135_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06789__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 total_design.keypad0.counter\[11\] vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11659__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10509_ net224 net2691 net483 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__mux2_1
X_14277_ net987 _01453_ net1083 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10563__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold619 total_design.core.regFile.register\[26\]\[1\] vssd1 vssd1 vccd1 vccd1 net1935
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11489_ net1603 _05621_ net149 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10790__C _05028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap349 _05819_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_4
XANTENNA__06613__Y _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13228_ clknet_leaf_168_clk _00695_ net1156 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06342__A _01915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13159_ clknet_leaf_176_clk _00626_ net1052 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_155_Left_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1308 total_design.core.regFile.register\[25\]\[5\] vssd1 vssd1 vccd1 vccd1 net2624
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1319 total_design.core.regFile.register\[26\]\[14\] vssd1 vssd1 vccd1 vccd1 net2635
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06961__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ _03227_ _03228_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__and2_2
XFILLER_0_109_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07651_ total_design.core.regFile.register\[21\]\[21\] net598 _03160_ _03161_ vssd1
+ vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_105_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06713__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09799__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06602_ total_design.core.regFile.register\[13\]\[1\] net666 net652 total_design.core.regFile.register\[7\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a22o_1
X_07582_ total_design.core.regFile.register\[25\]\[20\] net647 net581 total_design.core.regFile.register\[6\]\[20\]
+ _03095_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_157_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09321_ total_design.core.data_cpu_o\[12\] net755 _04560_ _04562_ _02024_ vssd1 vssd1
+ vccd1 vccd1 _04563_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_122_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06533_ net906 net888 _02028_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__nor3_1
XFILLER_0_125_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11470__A1 _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09252_ net250 net2757 net456 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__mux2_1
X_06464_ net744 net734 net732 vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08203_ total_design.core.data_mem.data_read_adr_reg\[17\] total_design.core.data_mem.data_read_adr_reg\[16\]
+ total_design.core.data_mem.data_read_adr_reg\[19\] total_design.core.data_mem.data_read_adr_reg\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__or4_1
XFILLER_0_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09183_ net706 _04429_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06395_ total_design.core.regFile.register\[23\]\[0\] net928 net912 net907 vssd1
+ vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout225_A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08134_ total_design.core.regFile.register\[5\]\[31\] net629 net563 total_design.core.regFile.register\[3\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__a22o_1
XANTENNA__07426__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11569__S net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11773__A2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ net750 _03559_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[29\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10473__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1134_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07016_ _02549_ _02551_ _02563_ net685 total_design.core.regFile.register\[0\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__o32a_4
XFILLER_0_141_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09266__C _04296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout594_A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07308__A_N _02818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ _04218_ _04219_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout761_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06952__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07918_ _03323_ _03327_ _03372_ _03371_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__a31o_1
X_08898_ net469 _02234_ _04151_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__o21ai_1
X_07849_ total_design.core.regFile.register\[16\]\[25\] net634 net598 total_design.core.regFile.register\[21\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__a22o_1
XANTENNA__06704__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860_ _05099_ _05104_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__xor2_2
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07370__X total_design.core.ctrl.imm_32\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09519_ _04391_ _04664_ _04687_ _04574_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__o22a_1
X_10791_ total_design.core.data_bus_o\[11\] total_design.core.data_bus_o\[13\] total_design.core.data_bus_o\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__or3_1
XANTENNA__10648__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12530_ net979 total_design.core.ctrl.instruction\[28\] net883 _01719_ vssd1 vssd1
+ vccd1 vccd1 _01567_ sky130_fd_sc_hd__a22o_1
XANTENNA__11461__A1 _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12461_ net1875 net165 net346 vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09406__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14200_ clknet_leaf_79_clk net1633 net1222 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
X_11412_ _01726_ _05030_ _05538_ _05608_ net513 vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_34_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09738__A _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ _01649_ _01650_ _01648_ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14131_ clknet_leaf_89_clk _01311_ net1260 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11479__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11343_ _05291_ _05459_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__or2_2
XANTENNA__10383__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08090__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14062_ clknet_leaf_101_clk _01242_ net1238 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[80\]
+ sky130_fd_sc_hd__dfrtp_1
X_11274_ _05524_ _05527_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__nand2b_1
XANTENNA__06162__A total_design.core.ctrl.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13013_ clknet_leaf_159_clk _00480_ net1142 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10225_ net2104 net391 vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07196__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ net244 net2585 net394 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5 total_design.core.data_mem.data_read_adr_reg\[9\] vssd1 vssd1 vccd1 vccd1 net1321
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10087_ net284 net2853 net402 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13915_ clknet_leaf_89_clk _01095_ net1263 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload3_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13846_ clknet_leaf_48_clk _01054_ net1098 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08817__A _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13777_ clknet_leaf_48_clk total_design.core.data_mem.stored_data_adr\[20\] net1102
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10558__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ _05217_ _05225_ _05221_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_100_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11452__A1 _05651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07656__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12728_ clknet_leaf_135_clk _00195_ net1189 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12659_ clknet_leaf_180_clk _00126_ net1042 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06180_ total_design.core.mem_ctrl.state\[1\] _01760_ vssd1 vssd1 vccd1 vccd1 total_design.core.mem_ctrl.next_state\[2\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_29_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold405 total_design.lcd_display.row_2\[15\] vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
X_14329_ clknet_leaf_38_clk _01490_ net1080 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10293__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold416 net85 vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold427 net93 vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold438 _01361_ vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 total_design.lcd_display.row_2\[9\] vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06503__C net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09870_ net206 net2321 net430 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__mux2_1
Xfanout907 _01963_ vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__buf_2
Xfanout918 net919 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 net930 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__buf_2
XANTENNA__07187__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _04071_ _04075_ _04060_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_146_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1105 total_design.core.regFile.register\[9\]\[31\] vssd1 vssd1 vccd1 vccd1 net2421
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1116 total_design.core.regFile.register\[26\]\[19\] vssd1 vssd1 vccd1 vccd1 net2432
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1127 total_design.core.regFile.register\[26\]\[6\] vssd1 vssd1 vccd1 vccd1 net2443
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ net308 total_design.core.data_mem.data_cpu_i\[18\] vssd1 vssd1 vccd1 vccd1
+ _04007_ sky130_fd_sc_hd__or2_1
Xhold1138 total_design.core.regFile.register\[9\]\[26\] vssd1 vssd1 vccd1 vccd1 net2454
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 total_design.core.regFile.register\[14\]\[30\] vssd1 vssd1 vccd1 vccd1 net2465
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07703_ total_design.core.regFile.register\[4\]\[22\] net621 net563 total_design.core.regFile.register\[3\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08683_ total_design.keypad0.counter\[16\] total_design.keypad0.counter\[17\] _03958_
+ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_124_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07634_ total_design.core.regFile.register\[11\]\[21\] net795 net777 total_design.core.regFile.register\[22\]\[21\]
+ _03145_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06698__A1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11424__Y _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11053__A1_N _05037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ total_design.core.regFile.register\[0\]\[19\] net875 _03066_ _03082_ vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[19\] sky130_fd_sc_hd__o22a_4
XANTENNA__10468__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout342_A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11153__A _05411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1084_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ _02742_ _04545_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_172_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11443__A1 _05609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06516_ total_design.core.regFile.register\[24\]\[0\] net747 net739 net725 vssd1
+ vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__and4_1
XANTENNA__07647__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06247__A _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07496_ total_design.core.regFile.register\[3\]\[18\] net865 net857 total_design.core.regFile.register\[18\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07111__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09235_ _04478_ _04479_ net702 vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11994__A2 _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06447_ net971 _01915_ _01917_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__or3_4
XANTENNA_fanout130_X net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1251_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09166_ _04191_ _04413_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__nand2_1
X_06378_ net926 net914 net910 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__and3_1
XANTENNA__06534__X _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08117_ total_design.core.regFile.register\[14\]\[31\] net862 _03605_ _03606_ _03608_
+ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08072__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09097_ _04344_ _04347_ net452 vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_43_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08181__B _03330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09992__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08048_ total_design.core.regFile.register\[2\]\[29\] net636 net620 total_design.core.regFile.register\[4\]\[29\]
+ _03533_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold950 total_design.core.regFile.register\[26\]\[27\] vssd1 vssd1 vccd1 vccd1 net2266
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout597_X net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold961 total_design.core.regFile.register\[8\]\[12\] vssd1 vssd1 vccd1 vccd1 net2277
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 total_design.core.regFile.register\[30\]\[7\] vssd1 vssd1 vccd1 vccd1 net2288
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 total_design.core.regFile.register\[2\]\[22\] vssd1 vssd1 vccd1 vccd1 net2299
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 total_design.core.regFile.register\[7\]\[8\] vssd1 vssd1 vccd1 vccd1 net2310
+ sky130_fd_sc_hd__dlygate4sd3_1
X_10010_ net191 net2154 net416 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__mux2_1
X_09999_ net229 net2740 net415 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08748__A1_N _03112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11961_ net709 _05822_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__nand2_2
XFILLER_0_98_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10912_ _05145_ _05169_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__xnor2_1
X_13700_ clknet_leaf_40_clk total_design.core.data_mem.stored_read_data\[7\] net1090
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[7\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07886__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ total_design.core.math.pc_val\[1\] _05771_ _05759_ vssd1 vssd1 vccd1 vccd1
+ _01445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07350__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13631_ clknet_leaf_61_clk total_design.core.data_mem.data_write_adr_i\[3\] net1129
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10843_ _05061_ _05086_ _05074_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_156_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10378__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11434__A1 _05679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07638__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13562_ clknet_leaf_125_clk _01029_ net1188 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10774_ net1266 total_design.core.data_bus_o\[27\] _05028_ vssd1 vssd1 vccd1 vccd1
+ _05033_ sky130_fd_sc_hd__and3_1
XFILLER_0_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08924__X _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12513_ net976 total_design.core.instr_mem.instruction_i\[20\] vssd1 vssd1 vccd1
+ vccd1 _01711_ sky130_fd_sc_hd__and2b_1
XFILLER_0_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13493_ clknet_leaf_158_clk _00960_ net1144 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_160_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_160_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08850__A2 total_design.core.ctrl.instruction\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11350__X _05609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12444_ net2059 net231 net347 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12375_ net991 _01634_ _01635_ _01636_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06163__Y _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14114_ clknet_leaf_87_clk _01294_ net1250 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11326_ _05580_ _05544_ _05559_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__or3b_1
XANTENNA__06613__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07810__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14045_ clknet_leaf_88_clk _01225_ net1249 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11257_ _05418_ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_128_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07169__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10208_ _04656_ net2324 net392 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11188_ _05439_ _05440_ _05443_ _05444_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_52_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13385__RESET_B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06620__A total_design.core.regFile.register\[29\]\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06916__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ net218 net2082 net398 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__mux2_1
XANTENNA__09315__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11672__S net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07877__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire310_A _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07341__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13829_ clknet_leaf_77_clk _01037_ net1216 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10288__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11425__A1 _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07629__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07350_ total_design.core.regFile.register\[30\]\[15\] net840 net788 total_design.core.regFile.register\[13\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06301_ _01808_ _01879_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__nor2_1
XANTENNA__10779__A3 total_design.core.data_bus_o\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07281_ total_design.core.regFile.register\[25\]\[14\] net650 net576 total_design.core.regFile.register\[24\]\[14\]
+ _02803_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_151_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_151_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09020_ _04271_ _04272_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__or2_1
X_06232_ net929 _01810_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11728__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06163_ net969 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__inv_2
XANTENNA__08054__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold202 total_design.core.data_mem.data_read_adr_reg2\[8\] vssd1 vssd1 vccd1 vccd1
+ net1518 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_117_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold213 total_design.lcd_display.row_1\[57\] vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold224 total_design.lcd_display.row_1\[96\] vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 total_design.lcd_display.row_1\[28\] vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold246 total_design.lcd_display.row_1\[95\] vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold257 total_design.lcd_display.row_1\[27\] vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 total_design.lcd_display.row_1\[40\] vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold279 total_design.lcd_display.row_1\[84\] vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ net280 total_design.core.regFile.register\[24\]\[4\] net422 vssd1 vssd1 vccd1
+ vccd1 _00235_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout704 net705 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout715 net716 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__buf_1
XANTENNA__12153__A2 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout726 net727 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_165_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09853_ net270 net2207 net431 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__mux2_1
Xfanout737 _02033_ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_165_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 _02030_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout292_A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06907__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout759 net762 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_8
X_08804_ total_design.core.data_mem.data_cpu_i\[1\] _02183_ total_design.core.data_mem.data_cpu_i\[2\]
+ net333 vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__a22o_1
X_09784_ net269 net2012 net439 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__mux2_1
X_06996_ _02496_ _02539_ _02536_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__o21a_1
XANTENNA__07580__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08735_ _02540_ _02589_ _03990_ _02118_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_1_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11582__S net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ total_design.lcd_display.cnt_500hz\[12\] _03944_ vssd1 vssd1 vccd1 vccd1
+ _03946_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07332__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07617_ total_design.core.regFile.register\[0\]\[20\] net873 _03123_ _03130_ vssd1
+ vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08597_ net1946 net339 net714 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[18\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__08176__B _03090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_X net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09987__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ total_design.core.regFile.register\[12\]\[19\] net773 net771 total_design.core.regFile.register\[28\]\[19\]
+ _03065_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06408__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout512_X net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07479_ total_design.core.regFile.register\[22\]\[18\] net674 net632 total_design.core.regFile.register\[16\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_142_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_142_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08832__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09218_ net312 _04142_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10490_ net169 net2000 net377 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_101_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09149_ total_design.core.math.pc_val\[5\] _04371_ vssd1 vssd1 vccd1 vccd1 _04398_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_134_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08045__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07399__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06424__B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12160_ total_design.core.math.pc_val\[2\] total_design.core.program_count.imm_val_reg\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11111_ net516 _05062_ _05365_ _05369_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__a31oi_1
X_12091_ total_design.lcd_display.row_2\[84\] _05818_ _05853_ total_design.lcd_display.row_2\[116\]
+ _05948_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_9_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10661__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold780 total_design.core.regFile.register\[7\]\[25\] vssd1 vssd1 vccd1 vccd1 net2096
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 total_design.core.regFile.register\[8\]\[4\] vssd1 vssd1 vccd1 vccd1 net2107
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11042_ _05212_ _05236_ _05238_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_110_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11104__B1 _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12993_ clknet_leaf_123_clk _00460_ net1167 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1480 total_design.core.regFile.register\[18\]\[28\] vssd1 vssd1 vccd1 vccd1 net2796
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09470__B net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1491 total_design.core.regFile.register\[25\]\[14\] vssd1 vssd1 vccd1 vccd1 net2807
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11944_ _05800_ net474 vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__nor2_4
XANTENNA__06439__X _02014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07323__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11875_ total_design.lcd_display.currentState\[5\] _05756_ net709 vssd1 vssd1 vccd1
+ vccd1 _01443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09897__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13614_ clknet_leaf_49_clk net1329 net1102 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10826_ _05079_ _05080_ _05083_ _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06318__C _01793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10757_ _01771_ _01773_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13545_ clknet_leaf_18_clk _01012_ net1048 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_133_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_133_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08814__B _02233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13476_ clknet_leaf_108_clk _00943_ net1223 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10688_ net171 net2090 net361 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12427_ _01681_ _01682_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09485__X _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ total_design.core.math.pc_val\[23\] net523 _01620_ _01621_ vssd1 vssd1 vccd1
+ vccd1 _01493_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11667__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11309_ _05566_ _05567_ _05564_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_77_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10571__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12289_ net993 _04653_ net895 vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12135__A2 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14028_ clknet_leaf_98_clk _01208_ net1246 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07547__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06850_ total_design.core.regFile.register\[22\]\[6\] net675 net595 total_design.core.regFile.register\[8\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07562__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_160_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06781_ net751 _02342_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[4\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_160_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06770__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08520_ _03856_ _03858_ _03870_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08451_ _03799_ _03804_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_69_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07402_ total_design.core.regFile.register\[27\]\[16\] net780 net768 total_design.core.regFile.register\[7\]\[16\]
+ _02928_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08382_ _03737_ _03738_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07333_ total_design.core.regFile.register\[9\]\[15\] net665 net622 total_design.core.regFile.register\[4\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_124_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08283__Y _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout138_A _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07264_ net970 _02696_ net967 vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09003_ net473 _02968_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__or2_1
X_06215_ total_design.core.instr_mem.instruction_adr_i\[25\] total_design.core.instr_mem.instruction_adr_stored\[25\]
+ net981 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07195_ total_design.core.regFile.register\[23\]\[12\] net810 net790 total_design.core.regFile.register\[24\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1047_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06146_ total_design.lcd_display.cnt_20ms\[4\] vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_167_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11582__A0 _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08740__A _03234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11577__S net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10481__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1214_A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12126__A2 _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout512 _01902_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ net201 net1975 net427 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__mux2_1
Xfanout523 net525 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__clkbuf_2
Xfanout534 net536 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_2
Xfanout545 _03672_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout674_A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout556 _04111_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09836_ net207 net2306 net434 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__mux2_1
Xfanout567 net568 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_4
Xfanout578 net580 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__buf_4
Xfanout589 net592 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07553__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ net212 net2248 net444 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__mux2_1
X_06979_ total_design.core.regFile.register\[16\]\[8\] net856 net778 total_design.core.regFile.register\[22\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__a22o_1
XANTENNA__06761__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout939_A _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08718_ total_design.keypad0.counter\[0\] total_design.keypad0.counter\[1\] total_design.keypad0.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__a21oi_1
X_09698_ net535 _04915_ _04921_ _04194_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__o22a_1
XFILLER_0_95_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08649_ total_design.lcd_display.cnt_500hz\[6\] _03933_ vssd1 vssd1 vccd1 vccd1 _03935_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_139_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06419__B total_design.core.ctrl.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11660_ _05627_ net1596 net130 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ net219 net2697 net365 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11591_ _05624_ net1639 net139 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10656__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_115_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13330_ clknet_leaf_137_clk _00797_ net1180 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10542_ net226 net2188 net376 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08018__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13261_ clknet_leaf_2_clk _00728_ net1014 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10473_ net239 net2277 net379 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12212_ total_design.core.math.pc_val\[7\] net528 _06058_ _06059_ vssd1 vssd1 vccd1
+ vccd1 _01477_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13192_ clknet_leaf_23_clk _00659_ net1057 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11573__A0 _05652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07777__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12143_ total_design.lcd_display.row_2\[71\] net349 _05839_ total_design.lcd_display.row_1\[63\]
+ _05997_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_92_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545__1267 vssd1 vssd1 vccd1 vccd1 _14545__1267/HI net1267 sky130_fd_sc_hd__conb_1
XFILLER_0_130_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10391__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12117__A2 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07792__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ total_design.lcd_display.row_1\[28\] _05838_ _05839_ total_design.lcd_display.row_1\[60\]
+ _03928_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11025_ _05272_ _05277_ _05273_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08809__B total_design.core.data_mem.data_cpu_i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12976_ clknet_leaf_185_clk _00443_ net1037 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11927_ total_design.keypad0.key_out\[7\] net529 net475 total_design.keypad0.key_out\[3\]
+ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11858_ _01724_ total_design.lcd_display.currentState\[1\] _05727_ _05729_ vssd1
+ vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_99_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09420__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10809_ _05065_ _05066_ _05063_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_64_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10566__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_106_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11789_ net1790 net954 net301 _01795_ vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13528_ clknet_leaf_133_clk _00995_ net1195 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_191_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13459_ clknet_leaf_177_clk _00926_ net1047 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__clkbuf_4
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11564__A0 _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09221__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07783__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ total_design.core.regFile.register\[23\]\[27\] net679 net617 total_design.core.regFile.register\[10\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06902_ total_design.core.regFile.register\[26\]\[7\] net644 net573 total_design.core.regFile.register\[24\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a22o_1
XANTENNA__06511__C net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07882_ total_design.core.regFile.register\[25\]\[26\] net843 net828 total_design.core.regFile.register\[1\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__a22o_1
XANTENNA__07535__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06833_ _02367_ _02389_ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09621_ _04508_ _04666_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__nand2_1
XANTENNA__06743__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ net197 net2530 net455 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__mux2_1
X_06764_ total_design.core.regFile.register\[4\]\[4\] net620 net562 total_design.core.regFile.register\[3\]\[4\]
+ _02325_ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08503_ _03834_ _03854_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__nand2_1
X_09483_ net903 _04717_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06695_ _02250_ _02253_ _02257_ _02261_ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__or4_1
X_08434_ _03787_ _03788_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_144_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06807__X _02367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08365_ net717 _03723_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[1\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_22_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10476__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout422_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10055__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07316_ total_design.core.ctrl.instruction\[15\] _02797_ vssd1 vssd1 vccd1 vccd1
+ _02847_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08296_ net1464 net941 _03682_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[5\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13488__RESET_B net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_159_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07247_ total_design.core.regFile.register\[12\]\[13\] _01980_ net776 total_design.core.regFile.register\[22\]\[13\]
+ _02774_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13417__RESET_B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12347__A2 _03234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07178_ _02701_ _02705_ _02706_ _02716_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout791_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09212__A2 _02515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout320 net321 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout331 net332 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_2
Xfanout342 net343 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_2
Xfanout353 _05018_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_4
Xfanout364 _05016_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__buf_4
Xfanout375 _05012_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_6
XANTENNA__09920__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 net387 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_8
X_09819_ net270 net2171 net436 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__mux2_1
Xfanout397 _04992_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06734__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12830_ clknet_leaf_180_clk _00297_ net1044 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12761_ clknet_leaf_188_clk _00228_ net1028 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14500_ clknet_leaf_36_clk _01567_ net1071 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[28\]
+ sky130_fd_sc_hd__dfrtp_4
X_11712_ net17 net934 net877 net2056 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__o22a_1
XFILLER_0_139_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12692_ clknet_leaf_141_clk _00159_ net1182 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11643_ _05628_ net1668 net136 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14431_ clknet_leaf_34_clk total_design.core.data_out_INSTR\[26\] net1067 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[26\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10386__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10046__A0 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11574_ _05636_ net1614 net144 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__mux2_1
X_14362_ clknet_leaf_10_clk _01503_ net1021 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_94_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
Xinput39 nrst vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_2
X_10525_ net163 net2076 net482 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__mux2_1
X_13313_ clknet_leaf_123_clk _00780_ net1167 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14293_ clknet_leaf_100_clk _01469_ net1231 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13244_ clknet_leaf_30_clk _00711_ net1060 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_131_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10456_ net172 net1993 net383 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ clknet_leaf_164_clk _00642_ net1164 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10387_ net187 net2275 net486 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12126_ total_design.lcd_display.row_2\[78\] _05806_ _05845_ total_design.lcd_display.row_2\[22\]
+ _05981_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06973__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ total_design.lcd_display.row_1\[27\] _05838_ _05843_ total_design.lcd_display.row_1\[123\]
+ _05824_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09911__A0 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ _05256_ _05261_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12510__A2 total_design.core.ctrl.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10788__C _05028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ clknet_leaf_181_clk _00426_ net1043 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11680__S net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10285__A0 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06480_ net741 net734 net733 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_103_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10296__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08150_ _03637_ _03638_ _03639_ _03640_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__or4_2
XFILLER_0_56_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09442__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07101_ net971 total_design.core.ctrl.instruction\[7\] _01918_ net888 net965 vssd1
+ vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__a32o_1
XFILLER_0_160_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08081_ total_design.core.regFile.register\[16\]\[30\] net856 _03570_ _03572_ _03574_
+ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07032_ total_design.core.regFile.register\[26\]\[9\] net871 net863 total_design.core.regFile.register\[14\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07756__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08846__C_N _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ net461 _04234_ _04235_ net326 _04233_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__o311a_1
XANTENNA__06964__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07934_ total_design.core.regFile.register\[22\]\[27\] net777 net766 total_design.core.regFile.register\[6\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__a22o_1
XANTENNA__07508__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07865_ _03364_ _03365_ _03366_ _03367_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__or4_1
XANTENNA__06716__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout372_A _05013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09604_ _03371_ net505 vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_127_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06816_ total_design.core.regFile.register\[9\]\[5\] net852 net807 total_design.core.regFile.register\[5\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__a22o_1
X_07796_ total_design.core.regFile.register\[0\]\[24\] net875 _03284_ _03301_ vssd1
+ vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_39_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06747_ total_design.core.regFile.register\[0\]\[4\] net873 _02303_ _02310_ vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[4\] sky130_fd_sc_hd__o22a_4
X_09535_ net465 _04729_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout160_X net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11590__S net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09130__A1 _02395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout637_A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09466_ _03038_ _04682_ _04700_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__o21ai_1
X_06678_ total_design.core.regFile.register\[2\]\[3\] net784 net760 total_design.core.regFile.register\[21\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__a22o_1
XANTENNA__06537__X _02111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08417_ net931 net932 vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09397_ net507 _04635_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout804_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10028__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08184__B _03467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09995__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ net1488 net939 _03708_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[31\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06416__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08279_ net1385 net557 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[29\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_46_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08912__B _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10310_ net233 net2394 net495 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07995__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11290_ _05505_ _05541_ _05545_ _05539_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09197__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07087__Y _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10241_ net242 net2855 net502 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10172_ net213 net2798 net394 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout961_X net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1104 net1105 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06955__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1115 net1116 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__clkbuf_4
Xfanout1126 net1128 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__clkbuf_4
Xfanout1137 net1144 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__buf_2
Xfanout150 _05682_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__buf_2
Xfanout1148 net1149 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout161 net162 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_2
Xfanout1159 net1162 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout172 net175 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_2
X_13931_ clknet_leaf_93_clk _01111_ net1255 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[77\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout183 net184 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_1
Xfanout194 net196 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__06707__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11700__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13862_ clknet_leaf_66_clk total_design.core.ctrl.imm_32\[1\] net1123 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07380__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12813_ clknet_leaf_0_clk _00280_ net1003 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13793_ clknet_leaf_113_clk total_design.core.data_mem.data_cpu_i\[2\] net1203 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10267__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10806__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12744_ clknet_leaf_169_clk _00211_ net1159 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07132__B1 _01986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06447__X _02022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09672__A2 _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12675_ clknet_leaf_5_clk _00142_ net1022 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14414_ clknet_leaf_35_clk total_design.core.data_out_INSTR\[9\] net1071 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ _05677_ net1705 net133 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14345_ clknet_leaf_44_clk _00032_ net1087 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11557_ _05635_ net1736 net142 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold609 _03966_ vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
X_10508_ net232 net2296 net481 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__mux2_1
X_14276_ net986 _01452_ net1087 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_11488_ net1568 _05477_ net152 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10439_ net241 net2676 net384 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__mux2_1
X_13227_ clknet_leaf_119_clk _00694_ net1171 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07199__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07738__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13158_ clknet_leaf_199_clk _00625_ net1001 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06946__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11675__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12109_ total_design.lcd_display.row_1\[101\] _05810_ _05852_ total_design.lcd_display.row_2\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__a22o_1
XANTENNA__07725__Y _03234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13089_ clknet_leaf_127_clk _00556_ net1170 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1309 total_design.core.regFile.register\[13\]\[24\] vssd1 vssd1 vccd1 vccd1 net2625
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10799__B _05028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07650_ total_design.core.regFile.register\[11\]\[21\] net613 net567 total_design.core.regFile.register\[12\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07371__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06601_ total_design.core.regFile.register\[4\]\[1\] net620 net562 total_design.core.regFile.register\[3\]\[1\]
+ _02156_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a221o_1
XANTENNA__07910__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07581_ total_design.core.regFile.register\[20\]\[20\] net670 net573 total_design.core.regFile.register\[24\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09320_ net904 _04561_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06532_ total_design.core.regFile.register\[0\]\[0\] net682 _02101_ _02105_ vssd1
+ vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_122_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1092 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09251_ net452 _04495_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06463_ _01924_ net901 _02018_ total_design.core.ctrl.instruction\[16\] total_design.core.ctrl.instruction\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__o311a_1
XFILLER_0_47_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08202_ total_design.core.data_mem.data_read_adr_reg\[21\] total_design.core.data_mem.data_read_adr_reg\[20\]
+ total_design.core.data_mem.data_read_adr_reg\[23\] total_design.core.data_mem.data_read_adr_reg\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__or4_1
XANTENNA__06517__B net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09182_ _02491_ _04428_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06394_ net927 net911 net907 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__and3_1
XFILLER_0_172_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11758__B1 _05037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08133_ total_design.core.regFile.register\[26\]\[31\] net645 net567 total_design.core.regFile.register\[12\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_170_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_6__f_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout218_A _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07977__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08064_ _03557_ _03558_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_31_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06533__A net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ total_design.core.regFile.register\[7\]\[9\] net654 _02553_ _02555_ _02562_
+ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_114_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_4__f_clk_X clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07729__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08926__A1 _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11585__S net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08966_ net473 _02868_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__or2_1
X_07917_ _03416_ _03417_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__or2_4
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ net334 _02286_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout754_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08179__B _03234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_95_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07848_ total_design.core.regFile.register\[30\]\[25\] net660 net602 total_design.core.regFile.register\[31\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_162_Right_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07901__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ total_design.core.regFile.register\[25\]\[24\] net843 net832 total_design.core.regFile.register\[31\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__a22o_1
XANTENNA__08907__B _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09518_ _04669_ _04750_ net328 vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__mux2_1
X_10790_ net34 total_design.core.data_bus_o\[12\] _05028_ vssd1 vssd1 vccd1 vccd1
+ _05049_ sky130_fd_sc_hd__and3_2
XANTENNA__07114__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08311__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11997__B1 _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _03040_ net701 _04684_ net533 vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06873__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12460_ net2644 net169 net344 vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09406__A2 _02918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11749__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11411_ net303 _05596_ _05653_ _05669_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__a31oi_4
X_12391_ _01648_ _01649_ _01650_ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__or3_1
XANTENNA__10664__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08642__B _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14130_ clknet_leaf_86_clk _01310_ net1248 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11342_ net302 _05472_ _05599_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_151_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06443__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11273_ _05522_ _05523_ _05531_ _05437_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_162_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14061_ clknet_leaf_91_clk _01241_ net1263 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_13012_ clknet_leaf_143_clk _00479_ net1175 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10224_ _04949_ net2776 net393 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06928__B1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11495__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09590__A1 total_design.core.ctrl.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10155_ net286 net1918 net394 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold6 total_design.core.data_mem.data_read_adr_reg\[1\] vssd1 vssd1 vccd1 vccd1 net1322
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10086_ _04116_ _04119_ _04972_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__or3_2
Xclkbuf_leaf_86_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10488__A0 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08145__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13914_ clknet_leaf_87_clk _01094_ net1247 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07353__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13845_ clknet_leaf_48_clk _01053_ net1102 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08817__B net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15__f_clk_X clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13776_ clknet_leaf_49_clk total_design.core.data_mem.stored_data_adr\[19\] net1103
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06618__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10988_ _05225_ _05246_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12727_ clknet_leaf_123_clk _00194_ net1166 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12658_ clknet_leaf_145_clk _00125_ net1179 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11609_ _05612_ net1737 net137 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__mux2_1
XANTENNA__10574__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12589_ clknet_leaf_2_clk _00056_ net1011 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10412__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_10_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14328_ clknet_leaf_39_clk _01489_ net1095 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06353__A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold406 total_design.lcd_display.row_2\[39\] vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold417 total_design.lcd_display.row_2\[21\] vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold428 net75 vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 total_design.lcd_display.row_2\[11\] vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14259_ clknet_leaf_95_clk _01438_ net1256 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.currentState\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06631__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06503__D net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06919__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout908 _01963_ vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_2
Xfanout919 _01927_ vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _04058_ _04059_ _04069_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_146_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07592__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_14__f_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold1106 total_design.core.regFile.register\[13\]\[19\] vssd1 vssd1 vccd1 vccd1 net2422
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 total_design.core.regFile.register\[13\]\[16\] vssd1 vssd1 vccd1 vccd1 net2433
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 total_design.core.regFile.register\[12\]\[3\] vssd1 vssd1 vccd1 vccd1 net2444
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ net308 total_design.core.data_mem.data_cpu_i\[18\] vssd1 vssd1 vccd1 vccd1
+ _04006_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_77_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1139 total_design.core.regFile.register\[25\]\[4\] vssd1 vssd1 vccd1 vccd1 net2455
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08136__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07702_ total_design.core.regFile.register\[30\]\[22\] net660 net602 total_design.core.regFile.register\[31\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08682_ total_design.keypad0.counter\[16\] _03958_ vssd1 vssd1 vccd1 vccd1 _03959_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07633_ total_design.core.regFile.register\[15\]\[21\] net847 net799 total_design.core.regFile.register\[29\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__a22o_1
XANTENNA__06698__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07564_ total_design.core.regFile.register\[25\]\[19\] net843 _03067_ _03070_ _03081_
+ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09097__B1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09303_ _02692_ _04544_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__and2_1
X_06515_ net745 net738 net724 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_172_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07495_ net308 vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__inv_2
XFILLER_0_174_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11721__X _05692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09234_ _02588_ _04477_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06446_ net971 _01918_ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__and2b_1
XFILLER_0_111_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09165_ _04411_ _04412_ net312 vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10484__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06377_ net920 net911 net946 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__and3_1
XANTENNA__06870__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12265__A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout502_A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08116_ total_design.core.regFile.register\[17\]\[31\] net820 _03607_ vssd1 vssd1
+ vccd1 vccd1 _03608_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09096_ net905 _04345_ _04346_ net752 _01751_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__o32a_2
XFILLER_0_114_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08047_ total_design.core.regFile.register\[10\]\[29\] net616 net573 total_design.core.regFile.register\[24\]\[29\]
+ _03541_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__a221o_1
XANTENNA__07280__C1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold940 total_design.core.regFile.register\[9\]\[2\] vssd1 vssd1 vccd1 vccd1 net2256
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 total_design.core.regFile.register\[13\]\[29\] vssd1 vssd1 vccd1 vccd1 net2267
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09574__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold962 total_design.core.regFile.register\[26\]\[25\] vssd1 vssd1 vccd1 vccd1 net2278
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold973 total_design.core.regFile.register\[6\]\[11\] vssd1 vssd1 vccd1 vccd1 net2289
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 total_design.core.regFile.register\[1\]\[9\] vssd1 vssd1 vccd1 vccd1 net2300
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 total_design.core.regFile.register\[20\]\[18\] vssd1 vssd1 vccd1 vccd1 net2311
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout969_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09572__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ net237 net2713 net415 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__mux2_1
XANTENNA__07583__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06202__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08949_ total_design.core.ctrl.instruction\[28\] total_design.core.ctrl.instruction\[29\]
+ total_design.core.ctrl.instruction\[31\] total_design.core.ctrl.instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_32_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08127__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ _05746_ _05754_ _05749_ _05742_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__or4b_1
XFILLER_0_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_174_Left_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10911_ _05104_ _05147_ _05148_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a21o_1
XANTENNA__06689__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ _05760_ _05768_ _05770_ _05764_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout924_X net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13630_ clknet_leaf_63_clk total_design.core.data_mem.data_write_adr_i\[2\] net1129
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12481__A_N net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10842_ _05100_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13561_ clknet_leaf_191_clk _01028_ net1029 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_55_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10773_ total_design.core.data_bus_o\[24\] net695 vssd1 vssd1 vccd1 vccd1 _05032_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07102__A3 _02022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12512_ net977 total_design.core.ctrl.instruction\[19\] net882 _01710_ vssd1 vssd1
+ vccd1 vccd1 _01558_ sky130_fd_sc_hd__a22o_1
X_13492_ clknet_leaf_143_clk _00959_ net1175 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12443_ net1943 net238 net346 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__mux2_1
XANTENNA__06861__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11198__A1 total_design.core.data_bus_o\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12374_ net991 _04840_ net895 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08940__X _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14113_ clknet_leaf_96_clk _01293_ net1253 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11325_ _05579_ _05583_ net294 vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06613__A2 total_design.core.data_mem.data_cpu_i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12147__B1 _05810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11256_ _05509_ _05510_ _05512_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__a21o_2
X_14044_ clknet_leaf_100_clk _01224_ net1229 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ _04635_ total_design.core.regFile.register\[16\]\[15\] net393 vssd1 vssd1
+ vccd1 vccd1 _00502_ sky130_fd_sc_hd__mux2_1
X_11187_ _05439_ _05440_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_52_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11370__A1 total_design.core.data_bus_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10138_ net214 net2838 net398 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_59_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08118__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10069_ net225 net2865 net408 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07326__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10569__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13828_ clknet_leaf_77_clk _01036_ net1216 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13759_ clknet_leaf_61_clk total_design.core.data_mem.stored_data_adr\[2\] net1130
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06300_ net964 _01878_ _01877_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10633__A0 _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10779__A4 total_design.core.data_bus_o\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07280_ total_design.core.regFile.register\[15\]\[14\] net607 _02812_ net686 vssd1
+ vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__a211o_1
XFILLER_0_127_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06231_ total_design.core.data_adr_o\[20\] _01809_ net961 vssd1 vssd1 vccd1 vccd1
+ _01810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06852__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08282__B net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06162_ total_design.core.ctrl.instruction\[19\] vssd1 vssd1 vccd1 vccd1 _01745_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_25_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold203 total_design.lcd_display.row_1\[5\] vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_117_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold214 total_design.lcd_display.row_1\[107\] vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06514__C net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06604__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold225 total_design.lcd_display.row_1\[9\] vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 total_design.lcd_display.row_1\[104\] vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__B1 _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold247 total_design.data_in_BUS\[12\] vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold258 total_design.lcd_display.row_1\[87\] vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 total_design.lcd_display.row_1\[127\] vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ net271 net2367 net423 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout705 _04204_ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__buf_2
XFILLER_0_1_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout716 _03905_ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07626__B _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ net276 net1909 net430 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__mux2_1
Xfanout727 _02045_ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__buf_2
Xfanout738 net739 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_165_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 net753 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__buf_2
X_08803_ total_design.core.data_mem.data_cpu_i\[0\] _02106_ total_design.core.data_mem.data_cpu_i\[1\]
+ _02183_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__o22a_1
X_09783_ net279 net2323 net440 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__mux2_1
X_06995_ total_design.core.ctrl.instruction\[21\] net889 _02028_ total_design.core.ctrl.instruction\[29\]
+ _02543_ vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[9\] sky130_fd_sc_hd__a221o_1
XANTENNA__09306__A1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ _02395_ _02442_ _02492_ _03989_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_1_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08738__A _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10479__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08665_ total_design.lcd_display.cnt_500hz\[12\] _03944_ vssd1 vssd1 vccd1 vccd1
+ _03945_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout452_A _04121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1194_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11164__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07616_ _03124_ _03126_ _03127_ _03129_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08596_ net1847 net338 net714 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[17\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_166_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12074__C1 _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07547_ total_design.core.regFile.register\[4\]\[19\] net814 net760 total_design.core.regFile.register\[21\]\[19\]
+ net692 vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07478_ total_design.core.regFile.register\[31\]\[18\] net601 net577 total_design.core.regFile.register\[27\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09217_ _04127_ _04462_ net316 vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06843__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06429_ total_design.core.regFile.register\[4\]\[0\] net758 _02000_ _01987_ _01981_
+ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout505_X net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09148_ total_design.core.math.pc_val\[5\] _04371_ vssd1 vssd1 vccd1 vccd1 _04397_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06424__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09079_ _04232_ _04234_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__or2_1
XANTENNA__12129__B1 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11110_ _01728_ _05362_ _05028_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__or3b_2
XANTENNA__08920__B _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12090_ total_design.lcd_display.row_2\[92\] _05837_ _05912_ _05947_ vssd1 vssd1
+ vccd1 vccd1 _05948_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_9_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold770 total_design.core.regFile.register\[21\]\[31\] vssd1 vssd1 vccd1 vccd1 net2086
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout874_X net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09735__C net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold781 total_design.core.regFile.register\[15\]\[23\] vssd1 vssd1 vccd1 vccd1 net2097
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ _05057_ _05261_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__nor2_1
Xhold792 total_design.core.regFile.register\[9\]\[27\] vssd1 vssd1 vccd1 vccd1 net2108
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09591__X _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07020__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11104__A1 total_design.core.data_bus_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12992_ clknet_leaf_1_clk _00459_ net1004 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1470 total_design.core.regFile.register\[18\]\[15\] vssd1 vssd1 vccd1 vccd1 net2786
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1481 total_design.core.regFile.register\[12\]\[28\] vssd1 vssd1 vccd1 vccd1 net2797
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11943_ _05750_ net531 vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__nand2_1
XANTENNA__10389__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1492 total_design.core.regFile.register\[1\]\[7\] vssd1 vssd1 vccd1 vccd1 net2808
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11874_ net531 vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__inv_2
XANTENNA__08935__X _04189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13613_ clknet_leaf_49_clk net1327 net1100 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10825_ net521 _05062_ _05074_ _05067_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__a31o_1
XFILLER_0_157_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07087__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13544_ clknet_leaf_171_clk _01011_ net1057 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12080__A2 _05804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10756_ total_design.core.regFile.register\[0\]\[31\] net355 vssd1 vssd1 vccd1 vccd1
+ _01030_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06455__X _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13475_ clknet_leaf_8_clk _00942_ net1018 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06174__Y _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10687_ net175 net2345 net363 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12426_ total_design.core.math.pc_val\[31\] net989 vssd1 vssd1 vccd1 vccd1 _01682_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12357_ net899 _03282_ net522 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__a21oi_1
XANTENNA_max_cap348_A _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11308_ _05554_ _05560_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12288_ _06113_ _06115_ _06116_ _06124_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__a211o_1
X_14027_ clknet_leaf_89_clk _01207_ net1259 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[109\]
+ sky130_fd_sc_hd__dfrtp_1
X_11239_ _05494_ _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_71_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07547__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07011__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11683__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06780_ _02315_ _02341_ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_160_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10299__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08450_ _03802_ _03803_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_69_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08845__X _04100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire306_X net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07401_ total_design.core.regFile.register\[3\]\[16\] net868 net836 total_design.core.regFile.register\[10\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__a22o_1
X_08381_ total_design.keypad0.key_out\[6\] total_design.keypad0.key_out\[4\] vssd1
+ vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__xor2_1
XFILLER_0_133_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07332_ total_design.core.regFile.register\[5\]\[15\] net630 net591 total_design.core.regFile.register\[1\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07078__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06365__X _01941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12071__A2 _05804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07263_ net970 net967 _02696_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__or3_1
XFILLER_0_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06825__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06214_ total_design.core.data_adr_o\[26\] _01792_ net962 vssd1 vssd1 vccd1 vccd1
+ _01793_ sky130_fd_sc_hd__mux2_1
XANTENNA__08747__A1_N _02918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09002_ _04253_ _04254_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09224__B1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07194_ total_design.core.regFile.register\[14\]\[12\] net863 net824 total_design.core.regFile.register\[19\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_115_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06145_ total_design.core.data_bus_o\[13\] vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08740__B _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07786__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07250__A2 _01932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06541__A _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09904_ net205 net2645 net426 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout502 net503 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__buf_6
XFILLER_0_111_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout513 net514 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_4
Xfanout524 net525 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_2
XFILLER_0_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout535 net536 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_4
Xfanout546 total_design.core.data_mem.next_write vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__buf_2
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout557 net558 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_2
X_09835_ net212 net1941 net436 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__mux2_1
XANTENNA__07002__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout568 _02092_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_8
Xfanout579 net580 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11593__S net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ net217 net2264 net442 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__mux2_1
X_06978_ total_design.core.regFile.register\[26\]\[8\] net871 net781 total_design.core.regFile.register\[27\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08717_ _03951_ _03978_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout834_A net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09697_ net295 _04578_ _04667_ _04575_ _04917_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__o221a_1
XANTENNA__08187__B _03602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09998__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10002__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08648_ _03933_ _03934_ net712 vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__and3b_1
XANTENNA__07710__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08579_ _03712_ _03906_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[0\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout622_X net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10610_ net215 net2741 net365 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07069__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12062__A2 _05826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11590_ _05635_ net1892 net138 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09463__B1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12840__RESET_B net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06816__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10541_ net234 net2420 net374 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13260_ clknet_leaf_170_clk _00727_ net1159 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10472_ net240 net2170 net377 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12211_ _02016_ _02492_ net526 vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_40_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10672__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13191_ clknet_leaf_18_clk _00658_ net1048 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07777__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12142_ total_design.lcd_display.row_1\[119\] _05814_ _05816_ total_design.lcd_display.row_1\[79\]
+ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__a22o_1
XANTENNA__06451__A total_design.core.ctrl.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07241__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12073_ net1601 net710 _05931_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__o21a_1
XANTENNA__07529__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11024_ _05275_ _05277_ _05272_ _05274_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06752__A1 total_design.core.ctrl.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12975_ clknet_leaf_147_clk _00442_ net1153 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06169__Y _01751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11926_ total_design.keypad0.key_out\[6\] net529 _05797_ total_design.keypad0.key_out\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__a22o_1
XANTENNA__07701__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11857_ total_design.lcd_display.currentState\[1\] _05742_ net709 vssd1 vssd1 vccd1
+ vccd1 _01439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10808_ _05065_ _05066_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__nand2_1
XANTENNA__06185__X _01766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11788_ net930 _01847_ _05698_ net956 net1542 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_64_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13527_ clknet_leaf_163_clk _00994_ net1165 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10739_ net2793 net354 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_136_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13458_ clknet_leaf_145_clk _00925_ net1179 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07480__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11678__S net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12409_ total_design.core.math.pc_val\[29\] net989 vssd1 vssd1 vccd1 vccd1 _01667_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_88_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10582__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__clkbuf_4
X_13389_ clknet_leaf_0_clk _00856_ net1005 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XANTENNA__07232__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07950_ total_design.core.regFile.register\[29\]\[27\] net657 net591 total_design.core.regFile.register\[1\]\[27\]
+ _03448_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_162_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06901_ total_design.core.regFile.register\[25\]\[7\] net647 net631 total_design.core.regFile.register\[5\]\[7\]
+ _02454_ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__a221o_1
X_07881_ total_design.core.regFile.register\[3\]\[26\] net867 net768 total_design.core.regFile.register\[7\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09620_ _03421_ net704 _04847_ net535 vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__a211o_1
X_06832_ _02389_ _02367_ vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07940__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ net452 _04782_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__nor2_1
X_06763_ total_design.core.regFile.register\[13\]\[4\] net666 net636 total_design.core.regFile.register\[2\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08502_ _03852_ _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__or2_1
X_09482_ _04715_ _04716_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__or2_1
X_06694_ _02242_ _02258_ _02259_ _02260_ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__or4_1
XANTENNA__07299__A2 _01947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08433_ _03785_ _03786_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout150_A _05682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09445__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08364_ total_design.data_in_BUS\[1\] net343 _03722_ vssd1 vssd1 vccd1 vccd1 _03723_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__12044__A2 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06536__A total_design.core.ctrl.imm_32\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07315_ total_design.core.ctrl.instruction\[15\] _02797_ vssd1 vssd1 vccd1 vccd1
+ _02846_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08295_ total_design.core.data_mem.data_write_adr_reg\[5\] net548 net541 total_design.core.data_mem.data_read_adr_reg\[5\]
+ net945 vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout415_A _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1157_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07246_ total_design.core.regFile.register\[1\]\[13\] net827 _02779_ _02780_ _02781_
+ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_171_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08751__A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11588__S net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10492__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07177_ total_design.core.regFile.register\[26\]\[12\] net646 _02715_ net688 vssd1
+ vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__a211o_1
XFILLER_0_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07223__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06271__A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout784_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout321 _02287_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout332 _02236_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_2
Xfanout343 _01905_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout572_X net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout354 _05018_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__buf_2
Xfanout365 net368 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_8
Xfanout376 _05012_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09381__C1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09818_ net278 net2549 net434 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__mux2_1
Xfanout387 net388 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_8
Xfanout398 _04990_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_6
X_09749_ net246 net1901 net443 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12760_ clknet_leaf_138_clk _00227_ net1184 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_6_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11711_ net16 net934 net877 net2148 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12691_ clknet_leaf_182_clk _00158_ net1041 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10667__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14430_ clknet_leaf_34_clk total_design.core.data_out_INSTR\[25\] net1067 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11642_ _05612_ net1618 net133 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12035__A2 _05804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14361_ clknet_leaf_30_clk _01502_ net1065 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11573_ _05652_ net1805 net143 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07998__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
X_13312_ clknet_leaf_1_clk _00779_ net1011 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_10524_ net166 net2105 net483 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14292_ clknet_leaf_94_clk _01468_ net1256 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07462__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11498__S net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13243_ clknet_leaf_149_clk _00710_ net1148 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10455_ net178 net2108 net383 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11546__A1 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13174_ clknet_leaf_155_clk _00641_ net1139 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10386_ net191 net2532 net486 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ total_design.lcd_display.row_1\[126\] _05843_ _05847_ total_design.lcd_display.row_2\[38\]
+ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12056_ total_design.lcd_display.row_2\[67\] net349 _05840_ total_design.lcd_display.row_1\[51\]
+ _05914_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _05257_ _05258_ _05265_ _05057_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__a211o_1
XANTENNA__07922__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ clknet_leaf_181_clk _00425_ net1044 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11909_ total_design.keypad0.next_rows\[1\] _05786_ _05785_ _05780_ vssd1 vssd1 vccd1
+ vccd1 _05787_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_138_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10577__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12889_ clknet_leaf_196_clk _00356_ net1009 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12026__A2 _05814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14559_ net1279 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_126_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11785__A1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07100_ _02641_ _02642_ net722 vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08080_ total_design.core.regFile.register\[13\]\[30\] net788 net769 total_design.core.regFile.register\[7\]\[30\]
+ _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07453__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07031_ total_design.core.regFile.register\[17\]\[9\] net821 net812 total_design.core.regFile.register\[23\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__a22o_1
XANTENNA__06661__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11537__A1 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08982_ net337 _02334_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07933_ total_design.core.regFile.register\[12\]\[27\] net773 net771 total_design.core.regFile.register\[28\]\[27\]
+ _03432_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout198_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09363__C1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ total_design.core.regFile.register\[13\]\[25\] net667 net637 total_design.core.regFile.register\[2\]\[25\]
+ _03351_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09603_ net322 _04750_ _04831_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_127_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06815_ total_design.core.regFile.register\[1\]\[5\] net829 _02373_ _02374_ vssd1
+ vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07795_ _03289_ _03291_ _03293_ _03300_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout365_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ _03228_ _04186_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_27_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06746_ _02305_ _02306_ _02307_ _02309_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__or4_1
XFILLER_0_64_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09130__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10487__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09465_ _03016_ _03035_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout153_X net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06677_ total_design.core.regFile.register\[26\]\[3\] net870 net807 total_design.core.regFile.register\[5\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08416_ net931 net932 vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12017__A2 _05834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07692__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ net904 _04633_ _04634_ _04632_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_4_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08347_ total_design.core.data_mem.data_write_adr_reg\[31\] net547 net539 total_design.core.data_mem.data_read_adr_reg\[31\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06416__D net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08278_ net1496 net558 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[28\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07444__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06652__B1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07229_ total_design.core.regFile.register\[7\]\[13\] net651 net650 total_design.core.regFile.register\[25\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11528__A1 _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07097__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10240_ net253 net2402 net500 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ net220 net2486 net396 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__mux2_1
Xfanout1105 net1135 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1116 net1121 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07825__A _03329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1127 net1128 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__buf_2
Xfanout140 _05685_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_2
Xfanout1138 net1144 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__clkbuf_4
Xfanout151 net152 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_4
Xfanout1149 net1154 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__clkbuf_2
Xfanout162 net164 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_2
X_13930_ clknet_leaf_85_clk _01110_ net1249 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_35_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout173 net174 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_2
Xfanout184 _04867_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07904__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout195 net196 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13861_ clknet_leaf_66_clk total_design.core.ctrl.imm_32\[0\] net1123 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_190_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12812_ clknet_leaf_174_clk _00279_ net1054 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13792_ clknet_leaf_113_clk total_design.core.data_mem.data_cpu_i\[1\] net1206 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11353__Y _05612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12743_ clknet_leaf_173_clk _00210_ net1054 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10397__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07683__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12674_ clknet_leaf_129_clk _00141_ net1197 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ clknet_leaf_38_clk total_design.core.data_out_INSTR\[8\] net1078 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[8\] sky130_fd_sc_hd__dfrtp_1
X_11625_ _05626_ net1673 net135 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14344_ clknet_leaf_46_clk _00031_ net1089 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11722__B1_N _05692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11556_ _05618_ net1856 net141 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__mux2_1
XANTENNA__07435__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__A _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10507_ net228 net1902 net480 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14275_ net986 _01451_ net1087 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_150_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07719__B _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11487_ _05674_ _05478_ _01855_ _05479_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__and4b_2
XANTENNA__11519__A1 _05630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ clknet_leaf_23_clk _00693_ net1057 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10438_ net253 net2846 net381 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12192__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ clknet_leaf_113_clk _00624_ net1203 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10369_ net266 net2859 net485 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_143_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12108_ _05958_ _05960_ _05962_ _05964_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13088_ clknet_leaf_194_clk _00555_ net1011 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08148__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12039_ total_design.lcd_display.row_2\[74\] _05806_ _05832_ total_design.lcd_display.row_2\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_158_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06600_ total_design.core.regFile.register\[25\]\[1\] net647 net570 total_design.core.regFile.register\[17\]\[1\]
+ _02158_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_105_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07580_ total_design.core.regFile.register\[9\]\[20\] net663 net632 total_design.core.regFile.register\[16\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06531_ _02096_ _02102_ _02103_ _02104_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_122_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09250_ _01756_ net752 _04494_ net905 _04493_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__o221a_2
XFILLER_0_47_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10100__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06462_ _01924_ net901 _02018_ _01744_ total_design.core.ctrl.instruction\[17\] vssd1
+ vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_174_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08201_ total_design.core.data_mem.state\[2\] _01749_ total_design.core.data_mem.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_174_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06882__B1 total_design.core.ctrl.imm_32\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06517__C net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09181_ _02390_ _02441_ _04403_ _04427_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06393_ _01739_ _01924_ net918 net908 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__and4_4
XFILLER_0_141_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09397__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08132_ _03599_ _03601_ _03598_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_170_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09820__A0 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07426__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06373__X _01949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06634__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08063_ _03507_ _03510_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__nor2_2
XFILLER_0_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07014_ total_design.core.regFile.register\[30\]\[9\] net661 _02559_ _02560_ _02561_
+ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_101_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12183__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11866__S net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08965_ net336 _02917_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout482_A _05011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08139__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ _03396_ _03415_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_87_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12486__A2 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08896_ net469 _02234_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__nor2_1
X_07847_ _03350_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[25\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__11454__X _05681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12613__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07778_ total_design.core.regFile.register\[12\]\[24\] net773 net771 total_design.core.regFile.register\[28\]\[24\]
+ _03283_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a221o_1
X_09517_ _04708_ _04749_ net468 vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06729_ total_design.core.regFile.register\[5\]\[4\] net806 net794 total_design.core.regFile.register\[11\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout535_X net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08311__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09448_ net701 _04683_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10010__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06873__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_96_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ _02892_ _04592_ _04616_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__nand3b_1
XANTENNA__08923__B net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11410_ net514 _05064_ _05459_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11749__B2 total_design.core.data_bus_o\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12390_ total_design.core.math.pc_val\[27\] net988 vssd1 vssd1 vccd1 vccd1 _01650_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06724__A _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06625__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11341_ _05459_ _05461_ _05466_ _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__o31a_1
XFILLER_0_90_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08090__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14060_ clknet_leaf_99_clk _01240_ net1229 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_11272_ _05524_ _05525_ _05527_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__a21o_2
XANTENNA__12174__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13011_ clknet_leaf_180_clk _00478_ net1041 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10223_ _04928_ net2419 net389 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__mux2_1
XANTENNA__10680__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07050__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10154_ _04115_ _04991_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_89_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 total_design.core.data_mem.data_read_adr_reg\[23\] vssd1 vssd1 vccd1 vccd1
+ net1323 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ net164 net2601 net408 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13913_ clknet_leaf_96_clk _01093_ net1254 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13844_ clknet_leaf_48_clk _01052_ net1103 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13775_ clknet_leaf_56_clk total_design.core.data_mem.stored_data_adr\[18\] net1115
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10987_ _05217_ _05223_ _05219_ _05218_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__o211ai_1
XANTENNA__06618__B _02188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12726_ clknet_leaf_153_clk _00193_ net1136 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07656__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06864__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12657_ clknet_leaf_150_clk _00124_ net1147 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11608_ _05609_ net1675 net139 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07408__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12588_ clknet_leaf_167_clk _00055_ net1155 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14327_ clknet_leaf_53_clk _01488_ net1095 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11539_ net1590 _05613_ net145 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08081__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold407 total_design.lcd_display.row_2\[96\] vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 total_design.lcd_display.row_2\[12\] vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14258_ clknet_leaf_43_clk net1415 net1082 vssd1 vssd1 vccd1 vccd1 wishbone.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
Xhold429 total_design.lcd_display.row_2\[75\] vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13209_ clknet_leaf_196_clk _00676_ net1009 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10590__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14189_ clknet_leaf_78_clk _01369_ net1217 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout909 net910 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07465__A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09581__A2 _03322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1107 total_design.core.regFile.register\[3\]\[23\] vssd1 vssd1 vccd1 vccd1 net2423
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08750_ _04000_ _04001_ _04002_ _04003_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__nand4_1
Xhold1118 total_design.core.regFile.register\[15\]\[24\] vssd1 vssd1 vccd1 vccd1 net2434
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 total_design.core.regFile.register\[3\]\[30\] vssd1 vssd1 vccd1 vccd1 net2445
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11676__A0 _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07701_ total_design.core.regFile.register\[9\]\[22\] net664 net598 total_design.core.regFile.register\[21\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__a22o_1
X_08681_ total_design.keypad0.counter\[15\] _03957_ vssd1 vssd1 vccd1 vccd1 _03958_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_124_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07632_ total_design.core.regFile.register\[16\]\[21\] net855 _03141_ _03142_ _03143_
+ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_36_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07895__A2 _03395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07563_ total_design.core.regFile.register\[24\]\[19\] net791 _03071_ _03074_ _03080_
+ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_165_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09302_ _02666_ _02687_ _04498_ _02637_ _04521_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06514_ total_design.core.regFile.register\[27\]\[0\] net748 net733 net725 vssd1
+ vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_172_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07494_ total_design.core.regFile.register\[0\]\[18\] net682 _03008_ _03014_ vssd1
+ vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__o22ai_2
XANTENNA__07647__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09233_ _02588_ _04477_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06855__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06445_ net896 _02019_ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__nand2_2
XFILLER_0_146_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07199__X total_design.core.data_mem.data_cpu_i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09164_ _04301_ _04304_ net324 vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__mux2_1
X_06376_ total_design.core.regFile.register\[9\]\[0\] net922 net915 net910 vssd1 vssd1
+ vccd1 vccd1 _01952_ sky130_fd_sc_hd__and4_1
XANTENNA__12265__B _02845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11600__A0 _05679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08115_ total_design.core.regFile.register\[19\]\[31\] net824 net765 total_design.core.regFile.register\[6\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09095_ total_design.core.math.pc_val\[2\] total_design.core.math.pc_val\[3\] vssd1
+ vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08072__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1237_A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08046_ total_design.core.regFile.register\[22\]\[29\] net674 net577 total_design.core.regFile.register\[27\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold930 total_design.core.regFile.register\[23\]\[24\] vssd1 vssd1 vccd1 vccd1 net2246
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11596__S net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold941 total_design.core.regFile.register\[7\]\[18\] vssd1 vssd1 vccd1 vccd1 net2257
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold952 total_design.core.regFile.register\[12\]\[2\] vssd1 vssd1 vccd1 vccd1 net2268
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold963 total_design.core.regFile.register\[8\]\[14\] vssd1 vssd1 vccd1 vccd1 net2279
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09574__B _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold974 total_design.core.regFile.register\[4\]\[28\] vssd1 vssd1 vccd1 vccd1 net2290
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold985 total_design.core.regFile.register\[27\]\[6\] vssd1 vssd1 vccd1 vccd1 net2301
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 total_design.core.regFile.register\[25\]\[0\] vssd1 vssd1 vccd1 vccd1 net2312
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07032__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ net241 net2178 net415 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10005__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ net285 net2711 net454 vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11667__A0 _05655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout652_X net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08879_ net334 _02770_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__nor2_1
XANTENNA__10800__Y _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ _05104_ _05147_ _05148_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09628__A2_N _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ _05769_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__inv_2
XANTENNA__07886__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10841_ _05061_ _05072_ _05085_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06438__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07099__B1 total_design.core.ctrl.instruction\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ clknet_leaf_135_clk _01027_ net1189 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[28\]
+ sky130_fd_sc_hd__dfrtp_2
X_10772_ total_design.core.data_bus_o\[26\] net695 vssd1 vssd1 vccd1 vccd1 _05031_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07638__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12511_ net977 total_design.core.instr_mem.instruction_i\[19\] vssd1 vssd1 vccd1
+ vccd1 _01710_ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06846__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13491_ clknet_leaf_180_clk _00958_ net1042 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10675__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12442_ net2041 net240 net344 vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11787__A2_N _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12373_ _01632_ _01633_ _01631_ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14112_ clknet_leaf_110_clk _01292_ net1226 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11324_ _05552_ _05582_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__nand2_1
XANTENNA__07271__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07810__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14043_ clknet_leaf_90_clk _01223_ net1261 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11255_ _05513_ _05509_ _05510_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_128_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10206_ _04614_ total_design.core.regFile.register\[16\]\[14\] net390 vssd1 vssd1
+ vccd1 vccd1 _00501_ sky130_fd_sc_hd__mux2_1
X_11186_ _05443_ _05444_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__nand2_1
XANTENNA__14441__RESET_B net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11370__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06620__C net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10137_ net221 net2567 net400 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11658__A0 _05626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10068_ net234 net2589 net409 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10330__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07877__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13827_ clknet_leaf_77_clk _01035_ net1130 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12083__B1 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13758_ clknet_leaf_59_clk total_design.core.data_mem.stored_data_adr\[1\] net1131
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07629__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08844__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ clknet_leaf_118_clk _00176_ net1160 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10585__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13689_ clknet_leaf_54_clk total_design.core.data_mem.data_read_adr_i\[29\] net1113
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06230_ total_design.core.instr_mem.instruction_adr_i\[20\] total_design.core.instr_mem.instruction_adr_stored\[20\]
+ net981 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10397__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06161_ total_design.core.ctrl.instruction\[18\] vssd1 vssd1 vccd1 vccd1 _01744_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_170_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08054__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08850__Y _04105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold204 total_design.lcd_display.row_1\[55\] vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold215 total_design.lcd_display.row_1\[43\] vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 net56 vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07801__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold237 total_design.lcd_display.row_1\[103\] vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold248 total_design.lcd_display.row_1\[7\] vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ net279 net2543 net423 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__mux2_1
Xhold259 total_design.lcd_display.row_1\[123\] vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout706 net708 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__clkbuf_4
Xfanout717 _03710_ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_2
XFILLER_0_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09851_ net244 net1935 net433 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__mux2_1
Xfanout728 net729 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_165_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 _02032_ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_2
XFILLER_0_147_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08802_ _04051_ _04054_ _04056_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__or3_1
X_09782_ net247 net2034 net438 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06994_ _02541_ _02542_ net722 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11649__A0 _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ _02188_ _02241_ _02292_ _02342_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08738__B _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout278_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09711__C1 _04105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ _03944_ net711 _03943_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__and3b_1
XFILLER_0_89_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11164__B _05184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07615_ total_design.core.regFile.register\[8\]\[20\] net802 _03128_ net691 vssd1
+ vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__a211o_1
X_08595_ total_design.data_in_BUS\[16\] net340 net714 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[16\]
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout445_A _04969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12074__B1 _05839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07546_ _03050_ _03063_ total_design.core.regFile.register\[0\]\[19\] net684 vssd1
+ vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_113_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08754__A _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10495__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08293__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07477_ total_design.core.regFile.register\[4\]\[18\] net620 net562 total_design.core.regFile.register\[3\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout612_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13810__D total_design.core.data_mem.data_cpu_i\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09216_ _04461_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__inv_2
X_06428_ _01739_ _01924_ net918 net908 vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__and4_1
XFILLER_0_91_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09147_ _04379_ _04394_ _04395_ net450 vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_32_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08045__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06359_ net951 net950 _01736_ total_design.core.ctrl.instruction\[21\] net952 vssd1
+ vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09078_ net969 _02289_ _02290_ net537 vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout981_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08029_ total_design.core.regFile.register\[17\]\[29\] net819 _01980_ total_design.core.regFile.register\[12\]\[29\]
+ _03524_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__a221o_1
Xhold760 total_design.core.regFile.register\[7\]\[31\] vssd1 vssd1 vccd1 vccd1 net2076
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold771 total_design.core.regFile.register\[26\]\[4\] vssd1 vssd1 vccd1 vccd1 net2087
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 total_design.core.regFile.register\[14\]\[25\] vssd1 vssd1 vccd1 vccd1 net2098
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11040_ _05212_ _05235_ _05238_ _05296_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__a31o_1
XANTENNA__06213__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold793 total_design.core.regFile.register\[13\]\[20\] vssd1 vssd1 vccd1 vccd1 net2109
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ clknet_leaf_155_clk _00458_ net1137 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11104__A2 _05049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1460 total_design.core.regFile.register\[16\]\[30\] vssd1 vssd1 vccd1 vccd1 net2776
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11942_ _05798_ _05803_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__nor2_4
XFILLER_0_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1471 total_design.core.regFile.register\[13\]\[12\] vssd1 vssd1 vccd1 vccd1 net2787
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1482 total_design.core.regFile.register\[17\]\[17\] vssd1 vssd1 vccd1 vccd1 net2798
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1493 total_design.core.regFile.register\[9\]\[12\] vssd1 vssd1 vccd1 vccd1 net2809
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06449__A total_design.core.ctrl.instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11873_ total_design.lcd_display.currentState\[5\] total_design.lcd_display.currentState\[3\]
+ _05723_ _05753_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__o31a_2
XFILLER_0_54_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13612_ clknet_leaf_56_clk net1350 net1115 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10824_ _05063_ _05067_ _05074_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__nand3b_1
XANTENNA__12065__B1 _05850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13543_ clknet_leaf_23_clk _01010_ net1055 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10755_ net2860 net356 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07492__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13474_ clknet_leaf_128_clk _00941_ net1194 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08951__X _04204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10686_ net177 net2360 net362 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12425_ _01674_ _01675_ _01672_ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08036__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07244__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ net991 _01617_ _01618_ _01619_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11307_ _05531_ _05562_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06190__Y _01770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12287_ _06124_ _06125_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14026_ clknet_leaf_86_clk _01206_ net1247 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[108\]
+ sky130_fd_sc_hd__dfrtp_1
X_11238_ _05493_ _05496_ _05490_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__a21o_1
XANTENNA__09062__A1_N total_design.core.data_cpu_o\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08744__B1 _01766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11169_ _05415_ _05417_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_143_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06770__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06522__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07400_ total_design.core.regFile.register\[18\]\[16\] net859 net792 total_design.core.regFile.register\[24\]\[16\]
+ _02926_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__a221o_1
X_08380_ _03735_ _03736_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__nand2_1
XANTENNA__12056__B1 _05840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold99_A total_design.bus_full vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07331_ total_design.core.regFile.register\[14\]\[15\] net626 net575 total_design.core.regFile.register\[24\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07262_ net751 _02796_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[13\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07483__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09001_ net335 _03112_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__or2_1
X_06213_ total_design.core.instr_mem.instruction_adr_i\[26\] total_design.core.instr_mem.instruction_adr_stored\[26\]
+ net981 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07193_ total_design.core.regFile.register\[12\]\[12\] net774 net772 total_design.core.regFile.register\[28\]\[12\]
+ _02731_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06144_ total_design.core.data_bus_o\[21\] vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_167_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08740__C _03330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09903_ net210 net2021 net427 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout503 _05003_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_4
Xfanout514 net515 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_2
Xfanout525 net528 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout395_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout536 _04106_ vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__buf_2
Xfanout547 total_design.core.data_mem.next_write vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_2
X_09834_ net218 net2544 net434 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__mux2_1
Xfanout558 net560 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_2
Xfanout569 _02091_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_8
X_09765_ net214 net2200 net442 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06977_ total_design.core.regFile.register\[12\]\[8\] net774 net772 total_design.core.regFile.register\[28\]\[8\]
+ _02527_ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout562_A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13805__D total_design.core.data_mem.data_cpu_i\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__06761__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ total_design.keypad0.counter\[3\] _03950_ vssd1 vssd1 vccd1 vccd1 _03978_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_69_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09696_ _04751_ _04920_ net320 vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__mux2_1
XANTENNA__07940__X total_design.core.data_mem.data_cpu_i\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08647_ total_design.lcd_display.cnt_500hz\[5\] _03931_ vssd1 vssd1 vccd1 vccd1 _03934_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_139_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout827_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08578_ _01775_ total_design.core.mem_ctrl.next_next_data_read total_design.core.mem_ctrl.next_next_fetch
+ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__or3b_2
XFILLER_0_7_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07529_ total_design.core.regFile.register\[19\]\[19\] net641 net583 total_design.core.regFile.register\[6\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10540_ net229 net2623 net374 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__mux2_1
XANTENNA__06208__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08018__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10471_ net255 net2687 net377 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_157_Right_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12210_ net994 _06055_ _06056_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__a31o_1
XANTENNA__07226__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13190_ clknet_leaf_198_clk _00657_ net1008 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09746__C total_design.core.ctrl.instruction\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout984_X net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ total_design.lcd_display.row_1\[39\] _05827_ _05840_ total_design.lcd_display.row_1\[55\]
+ _05995_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__a221o_1
XANTENNA__06434__D1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06451__B net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12072_ _05915_ _05918_ _05926_ _05930_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__or4_1
XFILLER_0_130_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold590 total_design.core.regFile.register\[6\]\[24\] vssd1 vssd1 vccd1 vccd1 net1906
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11023_ net351 _05055_ _05253_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_32_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12974_ clknet_leaf_189_clk _00441_ net1030 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08946__X _04200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1290 total_design.core.regFile.register\[26\]\[22\] vssd1 vssd1 vccd1 vccd1 net2606
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11925_ total_design.keypad0.key_out\[5\] net529 net475 total_design.keypad0.key_out\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12038__B1 _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ _05725_ _05735_ _05741_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_74_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ total_design.core.data_bus_o\[11\] total_design.core.data_bus_o\[13\] net698
+ net517 vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_99_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11787_ _01889_ _05693_ net953 net1689 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_28_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09454__A1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13526_ clknet_leaf_152_clk _00993_ net1138 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10738_ net2229 net353 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_41_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06345__C total_design.core.ctrl.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13457_ clknet_leaf_150_clk _00924_ net1147 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08009__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10669_ net254 net2701 net361 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12408_ _01656_ _01661_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__nand2_1
XANTENNA__07217__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ clknet_leaf_118_clk _00855_ net1160 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06642__A _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08560__C net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12339_ total_design.core.math.pc_val\[22\] total_design.core.program_count.imm_val_reg\[22\]
+ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__nand2_1
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XANTENNA__06976__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14009_ clknet_leaf_95_clk _01189_ net1254 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_06900_ total_design.core.regFile.register\[8\]\[7\] net596 net562 total_design.core.regFile.register\[3\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__a22o_1
X_07880_ total_design.core.regFile.register\[16\]\[26\] net855 net784 total_design.core.regFile.register\[2\]\[26\]
+ _03381_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_50_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07473__A total_design.core.ctrl.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_06831_ _02367_ _02389_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__or2_1
XANTENNA__06743__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ _02592_ _04776_ _04780_ _04781_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__and4_4
X_06762_ total_design.core.regFile.register\[10\]\[4\] net616 net585 total_design.core.regFile.register\[28\]\[4\]
+ _02323_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__a221o_1
XANTENNA__10103__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08501_ _03850_ _03851_ _03825_ _03830_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_108_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09481_ total_design.core.math.pc_val\[18\] _04676_ total_design.core.math.pc_val\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06693_ total_design.core.regFile.register\[13\]\[3\] net786 net763 total_design.core.regFile.register\[6\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__a22o_1
X_08432_ _03785_ _03786_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08363_ _01904_ _03720_ _03721_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__nor3_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout143_A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07314_ net751 _02845_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[14\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_22_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08294_ net1467 net941 _03681_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[4\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07245_ total_design.core.regFile.register\[14\]\[13\] net861 net850 total_design.core.regFile.register\[9\]\[13\]
+ _02773_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1052_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08751__B total_design.core.data_mem.data_cpu_i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07176_ total_design.core.regFile.register\[31\]\[12\] net603 net595 total_design.core.regFile.register\[8\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08956__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06271__B _01847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout777_A _01990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06982__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 net323 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_2
XANTENNA__10361__X _05007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout344 net347 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1105_X net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout355 _05018_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_4
Xfanout366 net368 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_8
Xfanout377 net380 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_6
X_09817_ net245 net1855 net435 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__mux2_1
Xfanout388 _05008_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout944_A _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07392__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout399 _04990_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout565_X net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06734__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ net285 net2101 net443 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09802__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ total_design.core.math.pc_val\[27\] total_design.core.math.pc_val\[28\] _04861_
+ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__and3_1
X_11710_ net15 net936 net879 net2839 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11491__A1 _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12690_ clknet_leaf_139_clk _00157_ net1184 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08645__C _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11641_ _05609_ net1777 net136 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14360_ clknet_leaf_45_clk _00029_ net1088 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07447__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11572_ _05613_ net1672 net141 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13311_ clknet_leaf_182_clk _00778_ net1040 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10523_ net169 net2220 net480 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__mux2_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_14291_ clknet_leaf_85_clk _01467_ net1251 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10683__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13242_ clknet_leaf_124_clk _00709_ net1188 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10454_ net182 net2454 net382 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08947__B1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13173_ clknet_leaf_166_clk _00640_ net1157 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10385_ net193 net2597 net484 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_107_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12124_ total_design.lcd_display.row_2\[62\] _05835_ _05978_ _05979_ vssd1 vssd1
+ vccd1 vccd1 _05980_ sky130_fd_sc_hd__a211o_1
XANTENNA__11367__X _05626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06973__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ total_design.lcd_display.row_1\[99\] _05810_ _05812_ total_design.lcd_display.row_1\[91\]
+ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__a22o_1
X_11006_ _05258_ _05260_ _05257_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09124__B1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ clknet_leaf_9_clk _00424_ net1019 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09675__B2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_116_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11908_ total_design.keypad0.next_rows\[3\] total_design.keypad0.next_rows\[2\] _03982_
+ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__and3_1
XANTENNA__11482__A1 _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07686__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ clknet_leaf_135_clk _00355_ net1186 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11839_ _05721_ _05722_ _05725_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14558_ net1278 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13509_ clknet_leaf_118_clk _00976_ net1171 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10593__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14489_ clknet_leaf_32_clk _01556_ net1063 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_130_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07030_ total_design.core.regFile.register\[12\]\[9\] _01994_ _01995_ total_design.core.regFile.register\[28\]\[9\]
+ _02577_ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07610__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ net470 _02286_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__nor2_1
X_07932_ total_design.core.regFile.register\[20\]\[27\] net816 net814 total_design.core.regFile.register\[4\]\[27\]
+ net692 vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__a221o_1
XANTENNA__07915__B _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12498__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07863_ total_design.core.regFile.register\[20\]\[25\] net671 net605 total_design.core.regFile.register\[15\]\[25\]
+ _03354_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__a221o_1
XANTENNA__06716__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06814_ total_design.core.regFile.register\[14\]\[5\] net863 net761 total_design.core.regFile.register\[21\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__a22o_1
X_09602_ net329 _04830_ _04196_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11156__C _05411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07794_ total_design.core.regFile.register\[19\]\[24\] net824 _03296_ _03298_ _03299_
+ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_127_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09533_ _03234_ net705 _04764_ net535 vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a211o_1
X_06745_ total_design.core.regFile.register\[23\]\[4\] net810 _02308_ net691 vssd1
+ vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout358_A _05017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11473__A1 _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ net217 net2662 net453 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06676_ total_design.core.regFile.register\[16\]\[3\] net924 vssd1 vssd1 vccd1 vccd1
+ _02243_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07141__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08415_ total_design.data_in_BUS\[5\] _01888_ net519 vssd1 vssd1 vccd1 vccd1 _03770_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09395_ total_design.core.ctrl.instruction\[15\] net886 net754 total_design.core.data_cpu_o\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout146_X net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08346_ net1501 net939 _03707_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[30\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07429__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08762__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11599__S net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08277_ net1381 net558 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[27\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_172_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14559__1279 vssd1 vssd1 vccd1 vccd1 _14559__1279/HI net1279 sky130_fd_sc_hd__conb_1
XFILLER_0_132_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07228_ total_design.core.regFile.register\[14\]\[13\] net624 net612 total_design.core.regFile.register\[11\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout894_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10008__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07159_ total_design.core.ctrl.instruction\[31\] _02028_ vssd1 vssd1 vccd1 vccd1
+ _02699_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1222_X net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07601__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10170_ net226 net2371 net396 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06955__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1106 net1108 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1117 net1120 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__clkbuf_4
Xfanout130 net131 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1128 net1133 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_3_6_0_clk_X clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout141 net142 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_4
Xfanout1139 net1144 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__clkbuf_2
Xfanout152 _05682_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06221__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout163 net164 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
Xfanout174 net175 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout185 net188 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06707__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout947_X net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11700__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 _04805_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_2
X_13860_ clknet_leaf_26_clk total_design.core.branch_ff net1107 vssd1 vssd1 vccd1
+ vccd1 total_design.core.program_count.ALU_out_reg sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07380__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12811_ clknet_leaf_119_clk _00278_ net1170 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10678__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13791_ clknet_leaf_113_clk total_design.core.data_mem.data_cpu_i\[0\] net1204 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11363__A _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12742_ clknet_leaf_197_clk _00209_ net1007 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07132__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12673_ clknet_leaf_121_clk _00140_ net1170 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_190_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_190_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_61_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _05624_ net1780 net135 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14412_ clknet_leaf_36_clk total_design.core.data_out_INSTR\[7\] net1084 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14343_ clknet_leaf_46_clk _00030_ net1088 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11555_ _05621_ net1514 net142 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__mux2_1
XANTENNA__08093__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10506_ net236 net2127 net481 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__mux2_1
XANTENNA__06643__A1 total_design.core.ctrl.instruction\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14274_ net987 _01450_ net1082 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07840__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06192__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11486_ net1562 _05630_ net156 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13225_ clknet_leaf_17_clk _00692_ net1046 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10437_ net252 net2295 net382 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ clknet_leaf_106_clk _00623_ net1234 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10368_ net273 net2499 net487 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__mux2_1
XANTENNA__06946__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12107_ total_design.lcd_display.row_1\[93\] _05812_ _05844_ total_design.lcd_display.row_2\[45\]
+ _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13087_ clknet_leaf_183_clk _00554_ net1039 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10299_ net268 net2325 net493 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12038_ total_design.lcd_display.row_1\[82\] _05815_ _05827_ total_design.lcd_display.row_1\[34\]
+ _05897_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08847__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07371__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10588__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13989_ clknet_leaf_92_clk _01169_ net1259 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06530_ total_design.core.regFile.register\[2\]\[0\] net636 _02067_ _02075_ _02057_
+ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_157_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11455__A1 _05477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07659__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06461_ net741 net738 net736 vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_174_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_181_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_181_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_174_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08200_ _03651_ _03654_ _03656_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__or3_2
XFILLER_0_91_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09180_ net311 _02438_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__nor2_1
XANTENNA__06882__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06392_ net926 net918 net908 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__and3_1
XFILLER_0_173_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08131_ _03622_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[31\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__08084__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09397__B _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08062_ _03553_ _03554_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__nand2_2
XFILLER_0_141_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07013_ total_design.core.regFile.register\[25\]\[9\] net649 net587 total_design.core.regFile.register\[28\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08964_ net289 _04216_ _04210_ _04208_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__o211a_1
XANTENNA__09275__A2_N net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1015_A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ _03396_ _03415_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__and2_1
X_08895_ _04145_ _04148_ net462 vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__mux2_1
X_07846_ total_design.core.regFile.register\[0\]\[25\] net875 _03336_ _03349_ vssd1
+ vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__o22ai_4
XANTENNA__07898__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__A _03253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10498__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ total_design.core.regFile.register\[20\]\[24\] net816 net814 total_design.core.regFile.register\[4\]\[24\]
+ net692 vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__a221o_1
XANTENNA__06570__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout642_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06728_ net751 _02292_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[3\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11446__A1 _05648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09516_ net472 _03178_ _04254_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07114__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14267__Q total_design.bus_full vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11997__A2 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09447_ _03038_ _04682_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06659_ total_design.core.regFile.register\[22\]\[2\] net674 net624 total_design.core.regFile.register\[14\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_172_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_172_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1172_X net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09378_ _04592_ _04616_ _02892_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_81_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11749__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ total_design.core.data_mem.data_write_adr_reg\[22\] net546 net538 total_design.core.data_mem.data_read_adr_reg\[22\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__a221o_1
XFILLER_0_163_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08075__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11340_ net294 _05597_ _05596_ _05594_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06216__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout897_X net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06443__C _01915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11271_ _05524_ _05525_ _05528_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13010_ clknet_leaf_145_clk _00477_ net1177 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12174__A2 _02292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10222_ _04909_ net2605 net392 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06928__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ _04119_ _04968_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_89_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input36_A gpio_in[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ net166 net1989 net408 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 total_design.core.data_mem.data_read_adr_reg\[22\] vssd1 vssd1 vccd1 vccd1
+ net1324 sky130_fd_sc_hd__dlygate4sd3_1
X_13912_ clknet_leaf_110_clk _01092_ net1227 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07353__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13843_ clknet_leaf_56_clk _01051_ net1115 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11437__A1 _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13774_ clknet_leaf_56_clk total_design.core.data_mem.stored_data_adr\[17\] net1115
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[17\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06187__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10986_ _05226_ _05231_ _05233_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__and3_1
XANTENNA__14177__Q net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12725_ clknet_leaf_158_clk _00192_ net1141 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_163_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_163_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_100_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12656_ clknet_leaf_186_clk _00123_ net1031 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11607_ _05636_ net1680 net139 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__mux2_1
XANTENNA__08066__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12587_ clknet_leaf_114_clk _00054_ net1202 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14326_ clknet_leaf_69_clk _01487_ net1109 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11538_ net1516 _05657_ net146 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold408 total_design.lcd_display.row_2\[88\] vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 total_design.lcd_display.row_1\[93\] vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11469_ net1606 _05655_ net153 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10724__X _05018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14257_ clknet_leaf_104_clk _01437_ net1234 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07746__A _03253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ clknet_leaf_133_clk _00675_ net1195 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14188_ clknet_leaf_79_clk _01368_ net1217 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06919__A2 _01951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13139_ clknet_leaf_179_clk _00606_ net1035 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07592__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09318__B1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1108 total_design.core.regFile.register\[2\]\[31\] vssd1 vssd1 vccd1 vccd1 net2424
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 total_design.core.regFile.register\[18\]\[21\] vssd1 vssd1 vccd1 vccd1 net2435
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07700_ total_design.core.regFile.register\[16\]\[22\] net634 net609 total_design.core.regFile.register\[18\]\[22\]
+ _03208_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08680_ total_design.keypad0.counter\[13\] total_design.keypad0.counter\[14\] _03956_
+ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__and3_1
XFILLER_0_174_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07344__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ total_design.core.regFile.register\[20\]\[21\] net816 net811 total_design.core.regFile.register\[23\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14558__1278 vssd1 vssd1 vccd1 vccd1 _14558__1278/HI net1278 sky130_fd_sc_hd__conb_1
XFILLER_0_36_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11428__A1 _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10111__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07562_ total_design.core.regFile.register\[22\]\[19\] net777 _03076_ _03078_ _03079_
+ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_48_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09301_ net241 net2707 net454 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__mux2_1
XANTENNA__09900__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06513_ net745 net732 net724 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07493_ _03010_ _03011_ _03012_ _03013_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_154_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_154_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09232_ _02539_ _04454_ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06444_ net973 net971 _01915_ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__or3_2
XFILLER_0_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09163_ _04305_ _04307_ net324 vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__mux2_1
XANTENNA__08057__B1 total_design.core.ctrl.imm_32\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06375_ net922 net914 net909 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__and3_4
XFILLER_0_161_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08114_ total_design.core.regFile.register\[23\]\[31\] net811 net807 total_design.core.regFile.register\[5\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09094_ total_design.core.math.pc_val\[2\] total_design.core.math.pc_val\[3\] vssd1
+ vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__and2_1
XANTENNA__07804__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08045_ total_design.core.regFile.register\[30\]\[29\] net659 net601 total_design.core.regFile.register\[31\]\[29\]
+ _03538_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold920 total_design.core.regFile.register\[28\]\[9\] vssd1 vssd1 vccd1 vccd1 net2236
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1132_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold931 total_design.core.regFile.register\[7\]\[7\] vssd1 vssd1 vccd1 vccd1 net2247
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 total_design.core.regFile.register\[13\]\[4\] vssd1 vssd1 vccd1 vccd1 net2258
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold953 total_design.core.regFile.register\[24\]\[16\] vssd1 vssd1 vccd1 vccd1 net2269
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 total_design.core.regFile.register\[26\]\[29\] vssd1 vssd1 vccd1 vccd1 net2280
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 total_design.core.regFile.register\[24\]\[31\] vssd1 vssd1 vccd1 vccd1 net2291
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 total_design.core.regFile.register\[10\]\[5\] vssd1 vssd1 vccd1 vccd1 net2302
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 total_design.core.regFile.register\[25\]\[28\] vssd1 vssd1 vccd1 vccd1 net2313
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09996_ net255 net2588 net414 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__mux2_1
X_14519__1291 vssd1 vssd1 vccd1 vccd1 net1291 _14519__1291/LO sky130_fd_sc_hd__conb_1
XANTENNA__07583__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ _04199_ _04200_ net506 vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__o21a_1
XANTENNA__06791__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout857_A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_X net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10810__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08878_ net470 _02718_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__nor2_1
XANTENNA__07335__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07391__A _02917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07829_ total_design.core.regFile.register\[8\]\[25\] net803 net765 total_design.core.regFile.register\[6\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout645_X net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ _05092_ _05096_ _05098_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__a21oi_4
XANTENNA__10021__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09810__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06438__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07099__A1 total_design.core.ctrl.instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10771_ net697 vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09493__C1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_145_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_145_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout812_X net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_142_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ net978 total_design.core.ctrl.instruction\[18\] net881 _01709_ vssd1 vssd1
+ vccd1 vccd1 _01557_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13490_ clknet_leaf_146_clk _00957_ net1177 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12441_ net2240 net253 net344 vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08048__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09796__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12395__A2 _03467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12372_ _01631_ _01632_ _01633_ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_157_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11323_ _05579_ _05581_ _05559_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__a21o_1
X_14111_ clknet_leaf_98_clk _01291_ net1242 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12147__A2 _05804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07566__A total_design.core.data_mem.data_cpu_i\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14042_ clknet_leaf_87_clk _01222_ net1250 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[124\]
+ sky130_fd_sc_hd__dfrtp_1
X_11254_ _05509_ _05512_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__nand2_1
XANTENNA__11359__Y _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14460__Q total_design.core.instr_mem.instruction_adr_i\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10205_ _04588_ net2795 net390 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11185_ _05356_ _05431_ _05435_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__nand3_1
XFILLER_0_66_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06620__D net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10136_ net226 net2786 net401 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__mux2_1
XANTENNA_input39_X net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10067_ net228 net1977 net406 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__mux2_1
XANTENNA__07326__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_5__f_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload1_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13826_ clknet_leaf_59_clk _01034_ net1131 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13757_ clknet_leaf_62_clk total_design.core.data_mem.stored_data_adr\[0\] net1131
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[0\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_136_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_136_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10969_ _05217_ _05225_ _05227_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12708_ clknet_leaf_128_clk _00175_ net1191 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13688_ clknet_leaf_56_clk total_design.core.data_mem.data_read_adr_i\[28\] net1113
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08563__C net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08039__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12639_ clknet_leaf_181_clk _00106_ net1043 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12386__A2 _03421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06160_ total_design.core.ctrl.instruction\[17\] vssd1 vssd1 vccd1 vccd1 _01743_
+ sky130_fd_sc_hd__inv_2
XANTENNA__11594__A0 _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08860__A total_design.core.ctrl.instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold205 net62 vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_117_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14309_ clknet_leaf_103_clk _00009_ net1237 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold216 total_design.lcd_display.row_1\[72\] vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 total_design.lcd_display.row_1\[60\] vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12138__A2 _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold238 total_design.lcd_display.row_1\[34\] vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold249 total_design.lcd_display.row_1\[118\] vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06470__C1 total_design.core.ctrl.instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout707 net708 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10106__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ net284 total_design.core.regFile.register\[26\]\[0\] net433 vssd1 vssd1 vccd1
+ vccd1 _00167_ sky130_fd_sc_hd__mux2_1
Xfanout718 net720 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_2
Xfanout729 _02044_ vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07565__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _04037_ _04040_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__or3_1
X_06993_ total_design.core.ctrl.instruction\[29\] _02493_ vssd1 vssd1 vccd1 vccd1
+ _02542_ sky130_fd_sc_hd__nand2_1
X_09781_ net285 total_design.core.regFile.register\[28\]\[0\] net441 vssd1 vssd1 vccd1
+ vccd1 _00103_ sky130_fd_sc_hd__mux2_1
XANTENNA__07970__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08732_ _03924_ _03925_ _03988_ vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.lcd_en
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_1_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12310__A2 _03040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08738__C _03040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ total_design.lcd_display.cnt_500hz\[11\] total_design.lcd_display.cnt_500hz\[10\]
+ _03941_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07614_ total_design.core.regFile.register\[22\]\[20\] net775 net763 total_design.core.regFile.register\[6\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__a22o_1
X_08594_ net1824 net338 net714 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[15\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_76_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07545_ _03052_ _03056_ _03062_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__nor3_1
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_127_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout438_A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07476_ total_design.core.regFile.register\[9\]\[18\] net663 net566 total_design.core.regFile.register\[12\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06427_ total_design.core.regFile.register\[7\]\[0\] net770 _01998_ _01957_ _01967_
+ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__a2111o_1
X_09215_ _04365_ _04460_ net326 vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout605_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09146_ net295 _04383_ _04388_ net298 vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__o22a_1
X_06358_ _01925_ _01928_ _01931_ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__or3_4
XFILLER_0_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11585__A0 _05630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09077_ _04159_ _04327_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06289_ total_design.core.data_adr_o\[5\] _01867_ net964 vssd1 vssd1 vccd1 vccd1
+ _01868_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1135_X net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10805__A total_design.core.data_bus_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12129__A2 _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08028_ total_design.core.regFile.register\[1\]\[29\] net827 net790 total_design.core.regFile.register\[24\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold750 total_design.core.regFile.register\[8\]\[6\] vssd1 vssd1 vccd1 vccd1 net2066
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout595_X net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold761 total_design.core.regFile.register\[25\]\[15\] vssd1 vssd1 vccd1 vccd1 net2077
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 total_design.core.regFile.register\[17\]\[20\] vssd1 vssd1 vccd1 vccd1 net2088
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold783 total_design.core.regFile.register\[29\]\[27\] vssd1 vssd1 vccd1 vccd1 net2099
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold794 total_design.core.regFile.register\[23\]\[21\] vssd1 vssd1 vccd1 vccd1 net2110
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10016__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09805__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06764__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ net177 net2159 net419 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ clknet_leaf_175_clk _00457_ net1053 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1450 total_design.core.regFile.register\[3\]\[24\] vssd1 vssd1 vccd1 vccd1 net2766
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 total_design.core.regFile.register\[21\]\[17\] vssd1 vssd1 vccd1 vccd1 net2777
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11941_ _05754_ _05802_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__or2_4
Xhold1472 total_design.core.regFile.register\[24\]\[8\] vssd1 vssd1 vccd1 vccd1 net2788
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1483 total_design.core.regFile.register\[10\]\[26\] vssd1 vssd1 vccd1 vccd1 net2799
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1494 total_design.core.regFile.register\[23\]\[31\] vssd1 vssd1 vccd1 vccd1 net2810
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11872_ total_design.lcd_display.currentState\[4\] _05754_ net709 vssd1 vssd1 vccd1
+ vccd1 _01442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13611_ clknet_leaf_58_clk net1341 net1118 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10823_ _05079_ _05080_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__or2_1
XANTENNA__10686__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_118_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13542_ clknet_leaf_195_clk _01009_ net1011 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_10754_ total_design.core.regFile.register\[0\]\[29\] net353 vssd1 vssd1 vccd1 vccd1
+ _01028_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08009__X _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14455__Q total_design.core.instr_mem.instruction_adr_i\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10685_ net182 net1959 net362 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__mux2_1
X_13473_ clknet_leaf_123_clk _00940_ net1167 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12424_ _04964_ _05757_ net527 vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_97_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06752__X total_design.core.ctrl.imm_32\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11576__A0 _05612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12355_ net991 _04801_ net895 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14557__1277 vssd1 vssd1 vccd1 vccd1 _14557__1277/HI net1277 sky130_fd_sc_hd__conb_1
XFILLER_0_26_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11306_ _05531_ _05562_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__nor2_1
X_12286_ _06113_ _06115_ _06116_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_147_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11237_ _05487_ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__nor2_1
X_14025_ clknet_leaf_96_clk _01205_ net1253 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_112_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10000__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07547__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11168_ net514 _05184_ _05424_ _05421_ _05420_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_143_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06755__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10119_ _04112_ _04119_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__nor2_1
X_11099_ net515 _05133_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__and2_2
XFILLER_0_117_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07180__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13809_ clknet_leaf_71_clk total_design.core.data_mem.data_cpu_i\[18\] net1205 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[18\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10596__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_109_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07330_ total_design.core.regFile.register\[15\]\[15\] net606 _02857_ _02858_ _02859_
+ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518__1290 vssd1 vssd1 vccd1 vccd1 net1290 _14518__1290/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_119_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07261_ _02751_ _02795_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_143_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09000_ net471 _03064_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__or2_1
X_06212_ total_design.core.data_adr_o\[30\] _01790_ net963 vssd1 vssd1 vccd1 vccd1
+ _01791_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07192_ total_design.core.regFile.register\[4\]\[12\] net815 net804 total_design.core.regFile.register\[8\]\[12\]
+ net693 vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__a221o_1
XANTENNA__11567__A0 _05679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06143_ total_design.core.data_bus_o\[16\] vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_167_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07786__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ net218 net2121 net429 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout504 net505 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__buf_2
XFILLER_0_10_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07538__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout526 net528 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_2
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09833_ net215 net2061 net434 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__mux2_1
Xfanout537 _04100_ vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_4
Xfanout548 total_design.core.data_mem.next_write vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_4
Xfanout559 net560 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_2
X_09764_ net223 net1940 net444 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__mux2_1
X_06976_ total_design.core.regFile.register\[19\]\[8\] net825 net815 total_design.core.regFile.register\[4\]\[8\]
+ net693 vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08715_ _03972_ _03975_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__nor2_1
X_09695_ _04830_ _04919_ net329 vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08646_ total_design.lcd_display.cnt_500hz\[5\] _03931_ vssd1 vssd1 vccd1 vccd1 _03933_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07171__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07710__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08577_ total_design.core.mem_ctrl.next_next_data_read total_design.core.mem_ctrl.next_next_fetch
+ _01774_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11102__D_N _01900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13821__D total_design.core.data_mem.data_cpu_i\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07528_ total_design.core.regFile.register\[14\]\[19\] net625 net571 total_design.core.regFile.register\[17\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07459_ total_design.core.regFile.register\[14\]\[17\] net864 net853 total_design.core.regFile.register\[28\]\[17\]
+ _02982_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1252_X net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_X net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10470_ net250 net2254 net379 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09129_ _02394_ _04376_ _04377_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_40_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09620__C1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ total_design.lcd_display.row_1\[7\] _05830_ _05994_ vssd1 vssd1 vccd1 vccd1
+ _05995_ sky130_fd_sc_hd__a21o_1
XANTENNA__07777__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06224__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10781__A1 total_design.core.data_bus_o\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06451__C _01915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__B1 total_design.core.ctrl.imm_32\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12071_ total_design.lcd_display.row_1\[67\] _05804_ _05847_ total_design.lcd_display.row_2\[35\]
+ _05929_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__a221o_1
XANTENNA__08785__A_N _02515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold580 total_design.core.regFile.register\[9\]\[13\] vssd1 vssd1 vccd1 vccd1 net1896
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07529__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold591 total_design.core.regFile.register\[25\]\[13\] vssd1 vssd1 vccd1 vccd1 net1907
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _05272_ _05278_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12522__A2 total_design.core.ctrl.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__06737__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12973_ clknet_leaf_6_clk _00440_ net1016 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1280 total_design.core.regFile.register\[26\]\[24\] vssd1 vssd1 vccd1 vccd1 net2596
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10297__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1291 total_design.core.regFile.register\[5\]\[11\] vssd1 vssd1 vccd1 vccd1 net2607
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11924_ total_design.keypad0.key_out\[4\] net530 net475 total_design.data_from_keypad\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__a22o_1
XANTENNA__06747__X total_design.core.data_mem.data_cpu_i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07162__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07701__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _05737_ _05739_ _05740_ total_design.lcd_display.currentState\[5\] vssd1
+ vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ total_design.core.data_bus_o\[11\] net699 _05059_ _05060_ net518 vssd1 vssd1
+ vccd1 vccd1 _05065_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11786_ net929 _01832_ _05694_ net953 net1505 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__a32o_1
XFILLER_0_144_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13525_ clknet_leaf_159_clk _00992_ net1143 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10737_ net2830 net353 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_136_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13456_ clknet_leaf_187_clk _00923_ net1031 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06482__X _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10668_ net251 net2141 net363 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ net900 _03559_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12210__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10599_ net272 net1913 net367 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__mux2_1
X_13387_ clknet_leaf_119_clk _00854_ net1171 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__clkbuf_4
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_140_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12338_ total_design.core.math.pc_val\[21\] net522 _01602_ _01603_ vssd1 vssd1 vccd1
+ vccd1 _01491_ sky130_fd_sc_hd__a22o_1
XANTENNA__12937__RESET_B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06976__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12269_ _06107_ _06108_ net993 vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__o21ai_1
X_14008_ clknet_leaf_74_clk _01188_ net1221 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09445__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06830_ _02108_ _02388_ _02347_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06761_ total_design.core.regFile.register\[29\]\[4\] net655 net640 total_design.core.regFile.register\[19\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a22o_1
X_08500_ _03825_ _03830_ _03850_ _03851_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__o211a_1
X_09480_ total_design.core.math.pc_val\[18\] total_design.core.math.pc_val\[19\] _04676_
+ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__and3_1
X_06692_ total_design.core.regFile.register\[3\]\[3\] net865 net767 total_design.core.regFile.register\[7\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__a22o_1
XANTENNA_wire311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09693__A2 _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08431_ total_design.keypad0.key_out\[10\] _03757_ _03755_ vssd1 vssd1 vccd1 vccd1
+ _03786_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06900__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08362_ total_design.keypad0.key_out\[1\] total_design.keypad0.key_out\[4\] _03719_
+ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08735__D _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07313_ _02843_ _02844_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__nand2_2
X_08293_ total_design.core.data_mem.data_write_adr_reg\[4\] net548 net541 total_design.core.data_mem.data_read_adr_reg\[4\]
+ net945 vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout136_A _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07244_ total_design.core.regFile.register\[11\]\[13\] net794 net758 total_design.core.regFile.register\[4\]\[13\]
+ _02772_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12201__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07175_ _02707_ _02709_ _02711_ _02713_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1045_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06967__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06431__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1212_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 _05700_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_2
Xfanout312 net315 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_2
XANTENNA__12504__A2 total_design.core.ctrl.instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout323 _02237_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_4
Xfanout334 net337 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_2
XANTENNA_fanout293_X net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06719__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout672_A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 net346 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_6
Xfanout356 _05018_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09381__A1 _02893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout367 net368 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_8
X_09816_ net286 net1893 net435 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__mux2_1
Xfanout378 net380 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_8
Xfanout389 net393 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07392__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ _04113_ _04116_ _04968_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__or3_4
XANTENNA__09669__C1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06959_ total_design.core.regFile.register\[14\]\[8\] net626 net622 total_design.core.regFile.register\[4\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout937_A _05688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09678_ _04895_ _04902_ _04903_ net450 vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14556__1276 vssd1 vssd1 vccd1 vccd1 _14556__1276/HI net1276 sky130_fd_sc_hd__conb_1
XFILLER_0_16_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08629_ net711 _03918_ _03919_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11640_ _05636_ net1652 net135 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__mux2_1
XANTENNA__06219__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_clk_X clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11571_ _05657_ net1772 net141 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08942__B _04193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07998__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13310_ clknet_leaf_180_clk _00777_ net1042 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10522_ net172 net1968 net482 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14290_ clknet_leaf_102_clk _01466_ net1238 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10453_ net185 net2390 net382 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__mux2_1
X_13241_ clknet_leaf_195_clk _00708_ net1010 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10203__A0 _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13172_ clknet_leaf_140_clk _00639_ net1183 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10384_ net199 net2230 net486 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__mux2_1
XANTENNA__06958__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12123_ total_design.lcd_display.row_2\[46\] _05844_ _05852_ total_design.lcd_display.row_2\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12054_ total_design.lcd_display.row_2\[27\] _05832_ _05845_ total_design.lcd_display.row_2\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__a22o_1
X_11005_ _05262_ _05263_ _05056_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10204__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06186__A1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07383__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout890 _02022_ vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__buf_2
XANTENNA__07922__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12956_ clknet_leaf_28_clk _00423_ net1073 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09675__A2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11907_ _05783_ _05784_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ clknet_leaf_161_clk _00354_ net1151 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ total_design.lcd_display.currentState\[3\] _05723_ _05724_ vssd1 vssd1 vccd1
+ vccd1 _05725_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14557_ net1277 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_155_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11769_ net1748 net956 net301 _01868_ vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_155_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10442__A0 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13508_ clknet_leaf_130_clk _00975_ net1198 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14488_ clknet_leaf_27_clk _01555_ net1074 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08571__C net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13439_ clknet_leaf_184_clk _00906_ net1039 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06661__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06949__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ _04211_ _04232_ net461 vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__or3b_1
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07931_ total_design.core.regFile.register\[5\]\[27\] net808 _03424_ _03429_ _03430_
+ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_48_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09363__A1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ total_design.core.regFile.register\[8\]\[25\] net594 net590 total_design.core.regFile.register\[1\]\[25\]
+ _03352_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__a221o_1
XANTENNA__10114__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08867__X _04121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07374__B1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09601_ net467 _04247_ _04250_ _04829_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__o31a_1
X_06813_ total_design.core.regFile.register\[8\]\[5\] net804 net785 total_design.core.regFile.register\[2\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07793_ total_design.core.regFile.register\[30\]\[24\] net839 net820 total_design.core.regFile.register\[17\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09532_ _04762_ _04763_ net707 vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__o21a_1
X_06744_ total_design.core.regFile.register\[31\]\[4\] net831 net786 total_design.core.regFile.register\[13\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07126__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06675_ total_design.core.regFile.register\[10\]\[3\] net836 net820 total_design.core.regFile.register\[17\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__a22o_1
X_09463_ _04695_ _04698_ net452 vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__a21oi_4
XANTENNA__06547__B net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08414_ net717 _03769_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[4\]
+ sky130_fd_sc_hd__nor2_1
X_09394_ total_design.core.math.pc_val\[15\] _04609_ vssd1 vssd1 vccd1 vccd1 _04633_
+ sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08345_ total_design.core.data_mem.data_write_adr_reg\[30\] net547 net539 total_design.core.data_mem.data_read_adr_reg\[30\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__a221o_1
XANTENNA__12422__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout420_A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1162_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout139_X net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08762__B _03322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06637__C1 _02190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08276_ net1491 net558 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[26\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06652__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07227_ total_design.core.regFile.register\[29\]\[13\] net658 _02760_ _02761_ _02762_
+ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07158_ _02696_ _02697_ net722 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08806__A1_N total_design.core.data_mem.data_cpu_i\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07089_ net551 net310 _02593_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout1215_X net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1107 net1108 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_2
Xfanout1118 net1120 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__clkbuf_4
Xfanout131 net132 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_4
Xfanout1129 net1133 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_98_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout142 _05684_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_4
Xfanout153 net154 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_4
XANTENNA__10024__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout164 _04967_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_35_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout175 _04910_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07904__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout186 net188 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout197 net200 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12810_ clknet_leaf_20_clk _00277_ net1050 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13790_ clknet_leaf_59_clk net549 net1127 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07117__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12110__B1 _05829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09657__A2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ clknet_leaf_119_clk _00208_ net1169 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12672_ clknet_leaf_1_clk _00139_ net1004 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14411_ clknet_leaf_41_clk total_design.core.data_out_INSTR\[6\] net1084 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _05635_ net1637 net134 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12413__A1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10694__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_133_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14342_ clknet_leaf_46_clk _00020_ net1088 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07569__A _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11554_ _05477_ net1723 net142 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10505_ net242 net2595 net481 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__mux2_1
X_14273_ net986 _01449_ net1082 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06192__B net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11485_ net1681 _05651_ net153 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13224_ clknet_leaf_173_clk _00691_ net1055 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10436_ net263 net2734 net383 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13155_ clknet_leaf_8_clk _00622_ net1020 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10367_ net258 net2080 net487 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__mux2_1
X_12106_ total_design.lcd_display.row_2\[21\] _05845_ _05847_ total_design.lcd_display.row_2\[37\]
+ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__a22o_1
X_10298_ net278 net2661 net493 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__mux2_1
X_13086_ clknet_leaf_175_clk _00553_ net1052 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_89_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08148__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12037_ total_design.lcd_display.row_1\[26\] _05838_ _05891_ _05895_ _05896_ vssd1
+ vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09950__C total_design.core.ctrl.instruction\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08847__B _04101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13988_ clknet_leaf_99_clk _01168_ net1241 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07108__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12101__B1 _05848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08305__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12939_ clknet_leaf_115_clk _00406_ net1202 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08856__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06367__B net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10663__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06460_ net742 net738 net736 vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_174_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06882__A2 total_design.core.data_mem.data_cpu_i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_84_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06391_ total_design.core.regFile.register\[17\]\[0\] net927 net948 net910 vssd1
+ vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_174_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08582__B net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08130_ total_design.core.regFile.register\[0\]\[31\] net875 _03621_ vssd1 vssd1
+ vccd1 vccd1 _03622_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_44_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08061_ _03553_ _03554_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06634__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10109__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07012_ total_design.core.regFile.register\[21\]\[9\] net599 net595 total_design.core.regFile.register\[8\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09033__A0 _02241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07766__X _03273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14555__1275 vssd1 vssd1 vccd1 vccd1 _14555__1275/HI net1275 sky130_fd_sc_hd__conb_1
XANTENNA__09584__B2 _04466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__A1 total_design.core.data_bus_o\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07595__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ net327 _04214_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08103__A _03595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08139__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07914_ _03399_ _03400_ _03414_ net684 total_design.core.regFile.register\[0\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__o32a_4
X_08894_ _04146_ _04147_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1008_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07845_ _03342_ _03344_ _03348_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout370_A _05013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__B _03273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09205__Y _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07776_ net749 _03282_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[23\]
+ sky130_fd_sc_hd__nor2_1
X_09515_ _03185_ net508 net448 _03182_ _04747_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__o221a_1
X_06727_ _02267_ _02291_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_149_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout635_A _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08311__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09446_ _02968_ _02989_ _02992_ _04638_ _04660_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__a221oi_2
X_06658_ _02219_ _02221_ _02223_ _02225_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__or4_1
XANTENNA__08773__A _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout802_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06873__A2 _01969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ _02818_ _02838_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__nand2_1
X_06589_ total_design.core.regFile.register\[31\]\[1\] net746 net732 net726 vssd1
+ vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__and4_1
XFILLER_0_163_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08328_ net1435 net938 _03698_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[21\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06625__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ net1386 net559 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[9\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_6_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09808__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11270_ _05524_ _05525_ _05528_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06580__X total_design.core.ctrl.imm_32\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10221_ _04889_ net391 _04999_ vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07586__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10152_ net163 net2593 net400 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__mux2_1
XANTENNA__07050__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10083_ net171 net2181 net406 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07338__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 total_design.core.data_mem.data_read_adr_reg\[14\] vssd1 vssd1 vccd1 vccd1
+ net1325 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13481__RESET_B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13911_ clknet_leaf_82_clk _01091_ net1220 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10689__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13842_ clknet_leaf_54_clk _01050_ net1109 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14458__Q total_design.core.instr_mem.instruction_adr_i\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13773_ clknet_leaf_56_clk total_design.core.data_mem.stored_data_adr\[16\] net1115
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[16\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12095__C1 _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ _05231_ _05233_ _05226_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06187__B total_design.core.instr_fetch vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08302__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12724_ clknet_leaf_141_clk _00191_ net1182 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07510__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12655_ clknet_leaf_161_clk _00122_ net1153 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06864__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11606_ _05652_ net1830 net140 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12586_ clknet_leaf_19_clk _00053_ net1050 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14325_ clknet_leaf_69_clk _01486_ net1109 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11537_ net1538 _05671_ net148 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold409 total_design.lcd_display.row_2\[19\] vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14256_ clknet_leaf_104_clk _01436_ net1234 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output97_A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ net1549 _05679_ net156 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13207_ clknet_leaf_164_clk _00674_ net1164 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10419_ net190 net2413 net386 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__mux2_1
X_14187_ clknet_leaf_79_clk _01367_ net1219 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11399_ _05361_ _05459_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__nand2_1
XANTENNA__07577__B1 total_design.core.ctrl.imm_32\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13569__RESET_B net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13138_ clknet_leaf_146_clk _00605_ net1178 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13069_ clknet_leaf_0_clk _00536_ net1006 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1109 total_design.core.regFile.register\[1\]\[18\] vssd1 vssd1 vccd1 vccd1 net2425
+ sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07329__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10599__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07630_ total_design.core.regFile.register\[8\]\[21\] net803 net765 total_design.core.regFile.register\[6\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07561_ total_design.core.regFile.register\[19\]\[19\] net824 net816 total_design.core.regFile.register\[20\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__a22o_1
X_09300_ net506 _04542_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__and2_1
X_06512_ total_design.core.regFile.register\[6\]\[0\] net743 net735 net731 vssd1 vssd1
+ vccd1 vccd1 _02086_ sky130_fd_sc_hd__and4_1
XFILLER_0_158_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07492_ total_design.core.regFile.register\[13\]\[18\] net666 net636 total_design.core.regFile.register\[2\]\[18\]
+ _02999_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__a221o_1
XANTENNA__07501__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09231_ _02515_ _02535_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06855__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06443_ net973 net971 _01915_ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__nor3_2
XFILLER_0_61_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06374_ net951 net950 total_design.core.ctrl.instruction\[20\] _01737_ net952 vssd1
+ vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__o2111a_2
X_09162_ _04408_ _04409_ net321 vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08113_ total_design.core.regFile.register\[12\]\[31\] net773 net771 total_design.core.regFile.register\[28\]\[31\]
+ _03604_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__a221o_1
XFILLER_0_161_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09093_ _04320_ _04334_ _04343_ net451 vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__a31o_1
XFILLER_0_142_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout216_A _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08044_ total_design.core.regFile.register\[9\]\[29\] net663 net566 total_design.core.regFile.register\[12\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__a22o_1
XANTENNA__07280__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold910 total_design.core.regFile.register\[11\]\[10\] vssd1 vssd1 vccd1 vccd1 net2226
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 total_design.core.regFile.register\[11\]\[1\] vssd1 vssd1 vccd1 vccd1 net2237
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold932 total_design.core.regFile.register\[29\]\[19\] vssd1 vssd1 vccd1 vccd1 net2248
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13992__RESET_B net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold943 total_design.core.regFile.register\[12\]\[12\] vssd1 vssd1 vccd1 vccd1 net2259
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 total_design.core.regFile.register\[4\]\[12\] vssd1 vssd1 vccd1 vccd1 net2270
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 total_design.core.regFile.register\[8\]\[18\] vssd1 vssd1 vccd1 vccd1 net2281
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 total_design.core.regFile.register\[30\]\[16\] vssd1 vssd1 vccd1 vccd1 net2292
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 total_design.core.regFile.register\[21\]\[29\] vssd1 vssd1 vccd1 vccd1 net2303
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 total_design.core.regFile.register\[29\]\[13\] vssd1 vssd1 vccd1 vccd1 net2314
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07032__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ net250 net2517 net417 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout585_A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08946_ total_design.core.math.pc_val\[0\] _02014_ net756 total_design.core.data_cpu_o\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__a22o_1
XANTENNA__08768__A total_design.core.data_mem.data_cpu_i\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07672__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06528__D1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ _04129_ _04130_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__nor2_1
XANTENNA__10810__B _05049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout752_A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07828_ total_design.core.regFile.register\[14\]\[25\] net862 net780 total_design.core.regFile.register\[27\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__a22o_1
XANTENNA__10302__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07740__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout540_X net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07759_ _03259_ _03261_ _03263_ _03265_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__or4_1
XFILLER_0_94_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10627__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout638_X net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10770_ net1266 _05028_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_143_Left_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09429_ _02337_ _04104_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06846__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12440_ net1988 net249 net346 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__mux2_1
XANTENNA__09245__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12371_ total_design.core.math.pc_val\[25\] net988 vssd1 vssd1 vccd1 vccd1 _01633_
+ sky130_fd_sc_hd__and2_1
X_14110_ clknet_leaf_101_clk _01290_ net1236 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11322_ _05552_ _05559_ _05544_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07847__A _03350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09538__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07271__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14041_ clknet_leaf_93_clk _01221_ net1253 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11253_ _05503_ _05511_ _05504_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_56_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07559__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_152_Left_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10204_ _04563_ net2463 net389 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07023__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ _05356_ _05438_ _05435_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_128_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10135_ net233 net2354 net399 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11107__A1 total_design.core.data_bus_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10066_ net237 net2828 net409 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__mux2_1
XANTENNA__10212__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07731__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13825_ clknet_leaf_59_clk _01033_ net1131 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11391__X _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_161_Left_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14554__1274 vssd1 vssd1 vccd1 vccd1 _14554__1274/HI net1274 sky130_fd_sc_hd__conb_1
XFILLER_0_156_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13756_ clknet_leaf_112_clk total_design.core.data_mem.stored_write_data\[31\] net1208
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[31\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__12083__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10968_ _05191_ _05197_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12707_ clknet_leaf_7_clk _00174_ net1016 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13687_ clknet_leaf_50_clk total_design.core.data_mem.data_read_adr_i\[27\] net1100
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[27\] sky130_fd_sc_hd__dfrtp_1
X_10899_ _05129_ _05138_ _05132_ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12638_ clknet_leaf_174_clk _00105_ net1053 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12569_ net1424 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14308_ clknet_leaf_103_clk _00008_ net1236 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold206 total_design.lcd_display.row_1\[81\] vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_117_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold217 total_design.lcd_display.row_1\[49\] vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold228 total_design.lcd_display.row_1\[82\] vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_170_Left_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14239_ clknet_leaf_57_clk _01419_ net1116 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold239 total_design.lcd_display.row_1\[92\] vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06380__B net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07014__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout719 net720 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__06222__A0 total_design.core.instr_mem.instruction_adr_i\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08800_ _04038_ _04039_ _04043_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__or3_1
X_09780_ _04113_ _04116_ _04118_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__or3_1
X_06992_ total_design.core.ctrl.instruction\[29\] _02493_ vssd1 vssd1 vccd1 vccd1
+ _02541_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07970__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ total_design.lcd_display.cnt_500hz\[3\] total_design.lcd_display.cnt_500hz\[2\]
+ total_design.lcd_display.cnt_500hz\[4\] vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11726__B _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09172__C1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10122__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08662_ total_design.lcd_display.cnt_500hz\[9\] total_design.lcd_display.cnt_500hz\[10\]
+ _03939_ total_design.lcd_display.cnt_500hz\[11\] vssd1 vssd1 vccd1 vccd1 _03943_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09911__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07613_ total_design.core.regFile.register\[18\]\[20\] net860 _01992_ total_design.core.regFile.register\[20\]\[20\]
+ _03116_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__a221o_1
X_08593_ net1857 net338 net714 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[14\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_89_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07544_ _03058_ _03060_ _03061_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__or3_1
XANTENNA__12074__A2 _05838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14191__RESET_B net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06828__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13730__Q total_design.core.data_bus_o\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07475_ total_design.core.ctrl.instruction\[30\] net885 net550 _02996_ vssd1 vssd1
+ vccd1 vccd1 total_design.core.ctrl.imm_32\[18\] sky130_fd_sc_hd__a211o_1
XFILLER_0_5_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1075_A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09214_ net460 _04143_ _04147_ _04459_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__o31a_1
XFILLER_0_146_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06426_ total_design.core.regFile.register\[16\]\[0\] net854 _01952_ _01965_ _01979_
+ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_107_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09145_ net289 _04391_ _04392_ _04393_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout500_A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06357_ net924 _01932_ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07789__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08770__B net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07667__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06288_ total_design.core.instr_mem.instruction_adr_i\[5\] total_design.core.instr_mem.instruction_adr_stored\[5\]
+ net984 vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__mux2_1
X_09076_ _04323_ _04326_ net319 vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08027_ _03516_ _03518_ _03520_ _03522_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__or4_1
Xhold740 total_design.data_in_BUS\[23\] vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 total_design.core.regFile.register\[16\]\[7\] vssd1 vssd1 vccd1 vccd1 net2067
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold762 total_design.core.regFile.register\[30\]\[30\] vssd1 vssd1 vccd1 vccd1 net2078
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 total_design.core.regFile.register\[26\]\[31\] vssd1 vssd1 vccd1 vccd1 net2089
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07005__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold784 total_design.core.regFile.register\[12\]\[11\] vssd1 vssd1 vccd1 vccd1 net2100
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold795 total_design.core.regFile.register\[29\]\[5\] vssd1 vssd1 vccd1 vccd1 net2111
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout588_X net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout967_A total_design.core.ctrl.instruction\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09978_ net181 net2754 net419 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07961__B1 total_design.core.ctrl.imm_32\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ _04179_ _04182_ net324 vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1440 total_design.core.regFile.register\[28\]\[24\] vssd1 vssd1 vccd1 vccd1 net2756
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1451 total_design.core.regFile.register\[5\]\[8\] vssd1 vssd1 vccd1 vccd1 net2767
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11940_ _05746_ _05749_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10032__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09702__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1462 total_design.core.regFile.register\[31\]\[21\] vssd1 vssd1 vccd1 vccd1 net2778
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1473 total_design.core.regFile.register\[16\]\[5\] vssd1 vssd1 vccd1 vccd1 net2789
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08010__B _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1484 total_design.core.regFile.register\[23\]\[20\] vssd1 vssd1 vccd1 vccd1 net2800
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1495 total_design.core.regFile.register\[23\]\[28\] vssd1 vssd1 vccd1 vccd1 net2811
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09821__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ _05750_ _05752_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__or2_4
XANTENNA__11652__A _05478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13610_ clknet_leaf_58_clk net1325 net1117 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10822_ _05079_ _05080_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__nor2_1
XANTENNA__12065__A2 _05834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13541_ clknet_leaf_116_clk _01008_ net1212 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10753_ total_design.core.regFile.register\[0\]\[28\] net355 vssd1 vssd1 vccd1 vccd1
+ _01027_ sky130_fd_sc_hd__and2_1
XANTENNA__06819__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ clknet_leaf_193_clk _00939_ net1012 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07492__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ net185 net2724 net362 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12423_ _01678_ _01679_ total_design.core.math.pc_val\[30\] net525 vssd1 vssd1 vccd1
+ vccd1 _01500_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_153_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14539__1311 vssd1 vssd1 vccd1 vccd1 net1311 _14539__1311/LO sky130_fd_sc_hd__conb_1
X_12354_ _01614_ _01616_ _01613_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07244__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10784__C1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11305_ _05548_ _05553_ _05563_ _05555_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__a31o_1
XANTENNA__11099__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12285_ _06122_ _06123_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10207__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14024_ clknet_leaf_111_clk _01204_ net1225 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[106\]
+ sky130_fd_sc_hd__dfrtp_1
X_11236_ _05389_ _05484_ _05482_ _05372_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06204__A0 total_design.core.instr_mem.instruction_adr_i\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11386__X _05645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07645__A2_N net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11167_ _05425_ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_143_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07952__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10118_ net162 net2603 net404 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11098_ _05356_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_160_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10049_ net170 net2303 net410 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__mux2_1
XANTENNA__09016__B _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11500__A1 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07704__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13808_ clknet_leaf_71_clk total_design.core.data_mem.data_cpu_i\[17\] net1206 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[17\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12056__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13739_ clknet_leaf_76_clk total_design.core.data_mem.stored_write_data\[14\] net1214
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07260_ _02794_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__inv_2
XANTENNA__07483__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06211_ total_design.core.instr_mem.instruction_adr_i\[30\] total_design.core.instr_mem.instruction_adr_stored\[30\]
+ net983 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06691__B1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07191_ total_design.core.regFile.register\[7\]\[12\] net769 _02729_ vssd1 vssd1
+ vccd1 vccd1 _02730_ sky130_fd_sc_hd__a21o_1
XANTENNA__09686__B _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11501__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06142_ total_design.core.mem_ctrl.state\[0\] vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10117__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09901_ net215 net2210 net426 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__mux2_1
XANTENNA__09906__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout505 _04187_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_4
Xfanout516 _01901_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout527 net528 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__buf_2
X_09832_ net221 net2731 net436 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_171_Right_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout538 _03676_ vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_2
XFILLER_0_10_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_141_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout549 total_design.core.data_mem.next_write vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07943__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ net224 net2412 net445 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__mux2_1
X_06975_ total_design.core.regFile.register\[5\]\[8\] net808 _02522_ _02524_ _02525_
+ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout283_A _04374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08714_ _03952_ _03977_ vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__and2b_1
XFILLER_0_174_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09694_ _04876_ _04918_ net468 vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08645_ _03931_ net712 _03928_ _03932_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout450_A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_156_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout548_A total_design.core.data_mem.next_write vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_166_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12047__A2 _05830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08576_ total_design.data_in_BUS\[31\] net340 net718 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[31\]
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07527_ total_design.core.regFile.register\[7\]\[19\] net653 net621 total_design.core.regFile.register\[4\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout715_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08120__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07458_ total_design.core.regFile.register\[25\]\[17\] net845 net794 total_design.core.regFile.register\[11\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06682__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06409_ total_design.core.regFile.register\[13\]\[0\] net923 net947 _01950_ vssd1
+ vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__and4_1
XFILLER_0_107_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07389_ _02902_ _02904_ _02914_ _02915_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09128_ _02394_ _04376_ net705 vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07226__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14291__Q net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10027__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09059_ net316 _04306_ _04310_ _04191_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06985__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10781__A2 total_design.core.data_bus_o\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09816__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12070_ total_design.lcd_display.row_2\[75\] _05806_ _05912_ _05928_ vssd1 vssd1
+ vccd1 vccd1 _05929_ sky130_fd_sc_hd__a211o_1
Xhold570 total_design.core.regFile.register\[15\]\[7\] vssd1 vssd1 vccd1 vccd1 net1886
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout872_X net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14553__1273 vssd1 vssd1 vccd1 vccd1 _14553__1273/HI net1273 sky130_fd_sc_hd__conb_1
Xhold581 total_design.core.regFile.register\[7\]\[1\] vssd1 vssd1 vccd1 vccd1 net1897
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 total_design.core.regFile.register\[16\]\[4\] vssd1 vssd1 vccd1 vccd1 net1908
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ _05272_ _05278_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12972_ clknet_leaf_166_clk _00439_ net1157 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1270 total_design.core.regFile.register\[6\]\[2\] vssd1 vssd1 vccd1 vccd1 net2586
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ _03981_ net999 net530 vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__a21oi_1
Xhold1281 total_design.core.regFile.register\[11\]\[23\] vssd1 vssd1 vccd1 vccd1 net2597
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1292 total_design.core.regFile.register\[11\]\[19\] vssd1 vssd1 vccd1 vccd1 net2608
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10697__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12038__A2 _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11854_ _05727_ _05734_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10805_ total_design.core.data_bus_o\[11\] net698 vssd1 vssd1 vccd1 vccd1 _05064_
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11785_ net929 _01816_ _05694_ net953 net1503 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08111__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13524_ clknet_leaf_143_clk _00991_ net1175 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10736_ net2667 net354 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13455_ clknet_leaf_161_clk _00922_ net1153 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ net262 net2819 net363 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__mux2_1
XANTENNA__11549__A1 _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12406_ total_design.core.math.pc_val\[28\] net524 _01663_ _01664_ vssd1 vssd1 vccd1
+ vccd1 _01498_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07217__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13386_ clknet_leaf_21_clk _00853_ net1050 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10598_ net258 net2035 net367 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10221__A1 _04889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__clkbuf_4
X_12337_ net899 _03187_ net522 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__a21oi_1
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_10_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12268_ _06107_ _06108_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14007_ clknet_leaf_83_clk _01187_ net1242 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11219_ _01903_ _05023_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_162_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12199_ _06045_ _06047_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__xor2_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07925__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08569__C net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06760_ total_design.core.regFile.register\[23\]\[4\] net678 net569 total_design.core.regFile.register\[17\]\[4\]
+ _02320_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__a221o_1
XANTENNA__09678__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06691_ total_design.core.regFile.register\[14\]\[3\] net861 net827 total_design.core.regFile.register\[1\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__a22o_1
X_08430_ _03783_ _03784_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__nand2_1
XANTENNA__10400__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08361_ total_design.keypad0.key_out\[4\] _03719_ total_design.keypad0.key_out\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08102__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11788__A1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07312_ _02791_ _02842_ _02841_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_22_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08292_ net1465 net940 _03680_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[3\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07243_ total_design.core.regFile.register\[19\]\[13\] net823 net763 total_design.core.regFile.register\[6\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__a22o_1
XANTENNA__07861__C1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout129_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07174_ total_design.core.regFile.register\[7\]\[12\] net652 net607 total_design.core.regFile.register\[15\]\[12\]
+ _02712_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12201__A2 _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08106__A _03595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06552__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1038_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_4
XANTENNA_fanout498_A _05004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7__f_clk_X clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout313 net315 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_2
Xfanout324 net325 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__buf_2
Xfanout335 net336 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_2
Xfanout346 net347 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_6
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout357 _05017_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_8
X_09815_ _04116_ _04971_ _04972_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__or3_4
Xfanout368 _05014_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_4
Xfanout379 net380 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout665_A _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout286_X net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ total_design.core.ctrl.instruction\[8\] net556 total_design.core.ctrl.instruction\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__nand3b_2
X_06958_ total_design.core.regFile.register\[9\]\[8\] net665 net635 total_design.core.regFile.register\[16\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14538__1310 vssd1 vssd1 vccd1 vccd1 net1310 _14538__1310/LO sky130_fd_sc_hd__conb_1
XFILLER_0_69_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09677_ _04552_ _04667_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__or2_1
X_06889_ _02028_ _02443_ total_design.core.ctrl.instruction\[27\] vssd1 vssd1 vccd1
+ vccd1 _02444_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout832_A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout453_X net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10310__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08628_ total_design.lcd_display.cnt_500hz\[1\] total_design.lcd_display.cnt_500hz\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__nand2_1
XANTENNA__07695__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout620_X net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08559_ net1857 net338 net718 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[14\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11570_ _05671_ net1676 net142 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__mux2_1
XANTENNA__07447__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10521_ net176 net2214 net482 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__mux2_1
XANTENNA__06655__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13240_ clknet_leaf_134_clk _00707_ net1195 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10452_ net191 net2576 net383 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08947__A2 _04200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13171_ clknet_leaf_178_clk _00638_ net1035 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10383_ net202 net2726 net486 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__mux2_1
X_12122_ total_design.lcd_display.row_2\[6\] _05850_ _05853_ total_design.lcd_display.row_2\[118\]
+ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07574__B _03090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12053_ _05803_ _05910_ _05911_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__and3_2
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07907__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ _05258_ _05260_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__and2b_1
XANTENNA__06186__A2 _01766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout880 _03906_ vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__buf_2
Xfanout891 _02022_ vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_clk sky130_fd_sc_hd__clkbuf_8
X_12955_ clknet_leaf_143_clk _00422_ net1173 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ total_design.keypad0.next_rows\[1\] _03983_ vssd1 vssd1 vccd1 vccd1 _05784_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_29_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07686__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12886_ clknet_leaf_153_clk _00353_ net1138 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ total_design.lcd_display.currentState\[5\] total_design.lcd_display.currentState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14556_ net1276 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11768_ net1625 net956 net301 _01861_ vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_155_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06934__A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06646__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10719_ net176 net2772 net359 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__mux2_1
X_13507_ clknet_leaf_7_clk _00974_ net1018 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14487_ clknet_leaf_32_clk _01554_ net1063 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_11699_ net3 net936 net879 net1882 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13438_ clknet_leaf_180_clk _00905_ net1044 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13369_ clknet_leaf_196_clk _00836_ net1009 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_max_cap349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07071__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07610__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07930_ total_design.core.regFile.register\[26\]\[27\] net871 net803 total_design.core.regFile.register\[8\]\[27\]
+ _03422_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__a221o_1
XANTENNA__09899__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12498__A2 total_design.core.ctrl.instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09363__A2 _04409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ total_design.core.regFile.register\[7\]\[25\] net653 _03363_ net687 vssd1
+ vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__a211o_1
X_09600_ net467 _04828_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__nand2_1
X_06812_ total_design.core.regFile.register\[29\]\[5\] net800 _02368_ _02371_ vssd1
+ vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__a211o_1
X_07792_ total_design.core.regFile.register\[10\]\[24\] net835 _03297_ vssd1 vssd1
+ vccd1 vccd1 _03298_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09531_ _03230_ _04744_ _04761_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__nor3_1
XANTENNA__09044__X _04296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06743_ total_design.core.regFile.register\[14\]\[4\] net861 net798 total_design.core.regFile.register\[29\]\[4\]
+ _02294_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10130__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09462_ net903 _04696_ _04697_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__o21ba_1
X_06674_ net751 _02241_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[2\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08413_ _03766_ _03767_ _03750_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06547__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09393_ _04620_ _04630_ _04631_ net449 vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__a31o_1
XFILLER_0_164_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout246_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14552__1272 vssd1 vssd1 vccd1 vccd1 _14552__1272/HI net1272 sky130_fd_sc_hd__conb_1
XFILLER_0_164_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08344_ net1462 net938 _03706_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[29\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07429__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12422__A2 _03602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11630__A0 _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06637__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08275_ net1401 net558 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[25\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_7_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1155_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07226_ total_design.core.regFile.register\[8\]\[13\] net593 net577 total_design.core.regFile.register\[27\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07157_ total_design.core.ctrl.instruction\[12\] _02641_ vssd1 vssd1 vccd1 vccd1
+ _02697_ sky130_fd_sc_hd__nand2_1
XANTENNA__07062__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07088_ net310 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[10\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__07601__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1108 net1135 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__buf_2
XANTENNA__10305__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1119 net1120 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__clkbuf_2
Xfanout132 _05687_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_2
Xclkbuf_4_1__f_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xfanout143 net144 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_4
Xfanout154 _05681_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout570_X net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout165 _04950_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_2
Xfanout176 net179 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout187 net188 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_2
Xfanout198 net200 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_87_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09729_ _03645_ _04951_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10040__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12740_ clknet_leaf_130_clk _00207_ net1198 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10121__A0 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08865__A1 total_design.core.ctrl.instruction\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12671_ clknet_leaf_155_clk _00138_ net1137 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14410_ clknet_leaf_41_clk total_design.core.data_out_INSTR\[5\] net1090 vssd1 vssd1
+ vccd1 vccd1 total_design.core.instr_mem.instruction_i\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11622_ _05618_ net1775 net133 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ clknet_leaf_44_clk _00004_ net1087 vssd1 vssd1 vccd1 vccd1 total_design.key_confirm
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06628__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11553_ _05478_ _05479_ _05674_ _05675_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_133_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08093__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06473__B _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10504_ net255 net2702 net480 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__mux2_1
X_14272_ net986 _01448_ net1085 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_52_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11484_ net1735 _05650_ net156 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07840__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06192__C total_design.core.instr_fetch vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13223_ clknet_leaf_176_clk _00690_ net1058 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10435_ net266 net2232 net381 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__mux2_1
XANTENNA__10188__A0 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_950 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13154_ clknet_leaf_129_clk _00621_ net1197 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10366_ net283 net2102 net484 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12105_ total_design.lcd_display.row_2\[69\] net349 _05850_ total_design.lcd_display.row_2\[5\]
+ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_29_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06800__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13085_ clknet_leaf_15_clk _00552_ net1025 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10297_ net246 net1853 net492 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__mux2_1
XANTENNA__07872__X _03375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12036_ total_design.lcd_display.row_1\[74\] _05816_ _05826_ total_design.lcd_display.row_1\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__a22o_1
XANTENNA__12172__C_N net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06488__X _02062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09305__A _02746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08305__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13987_ clknet_leaf_92_clk _01167_ net1253 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07659__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12938_ clknet_leaf_23_clk _00405_ net1057 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08856__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_38_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06367__C net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06867__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12869_ clknet_leaf_117_clk _00336_ net1171 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06390_ net925 net948 net909 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_174_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11612__A0 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14539_ net1311 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XANTENNA__08084__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07292__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08060_ _03554_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07831__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07011_ total_design.core.regFile.register\[20\]\[9\] net672 _02556_ _02558_ net688
+ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12992__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07495__A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11391__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10125__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ _04214_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__inv_2
X_07913_ _03402_ _03404_ _03406_ _03413_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__or4_1
XANTENNA__09914__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11679__A0 _05645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08893_ net334 _02367_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07844_ total_design.core.regFile.register\[15\]\[25\] net847 _03345_ _03347_ vssd1
+ vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__a211o_1
XANTENNA__06398__X _01974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07898__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07775_ _03280_ _03281_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__nand2_4
XANTENNA__13733__Q total_design.core.data_bus_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout363_A net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06570__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09514_ _03183_ net505 vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_56_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06726_ _02289_ _02290_ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__and2_2
XFILLER_0_66_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ net215 net2205 net453 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__mux2_1
XANTENNA__06858__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06657_ total_design.core.regFile.register\[10\]\[2\] net618 net585 total_design.core.regFile.register\[28\]\[2\]
+ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout151_X net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout628_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08773__B _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09376_ net232 net2349 net454 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06588_ total_design.core.regFile.register\[11\]\[1\] net740 net732 net723 vssd1
+ vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__and4_1
XFILLER_0_164_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11603__A0 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08327_ total_design.core.data_mem.data_write_adr_reg\[21\] net546 net538 total_design.core.data_mem.data_read_adr_reg\[21\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__a221o_1
XFILLER_0_163_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08075__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06293__B _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07283__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08258_ net1390 net559 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[8\]
+ sky130_fd_sc_hd__and2_1
X_07209_ net751 _02746_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[12\]
+ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_65_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07676__Y _03187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08189_ net1478 _01749_ net982 vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a21oi_1
X_10220_ net2640 net391 vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10151_ net165 net2106 net401 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10035__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09824__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10082_ net172 net2386 net408 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__mux2_1
Xwire1000 _05775_ vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910_ clknet_leaf_101_clk _01090_ net1237 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07889__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ clknet_leaf_56_clk _01049_ net1115 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13772_ clknet_leaf_58_clk total_design.core.data_mem.stored_data_adr\[15\] net1118
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[15\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12095__B1 _05839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10984_ _05208_ _05210_ _05240_ _05242_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__nand4_1
XFILLER_0_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06849__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12723_ clknet_leaf_179_clk _00190_ net1042 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11390__A _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ clknet_leaf_187_clk _00121_ net1028 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11605_ _05613_ net1928 net137 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12585_ clknet_leaf_17_clk _00052_ net1046 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08066__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11536_ net1581 _05680_ net147 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__mux2_1
X_14324_ clknet_leaf_69_clk _01485_ net1107 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07274__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07813__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11389__X _05648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14255_ clknet_leaf_104_clk _01435_ net1234 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11467_ net1607 _05632_ net154 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13206_ clknet_leaf_153_clk _00673_ net1138 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07026__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10418_ net195 net2428 net385 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14186_ clknet_leaf_79_clk _01366_ net1218 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfrtp_1
X_11398_ net513 _05608_ _05656_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__nand3_4
XFILLER_0_110_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13137_ clknet_leaf_150_clk _00604_ net1147 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10349_ net207 net2070 net488 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__mux2_1
XANTENNA__09019__B _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14551__1271 vssd1 vssd1 vccd1 vccd1 _14551__1271/HI net1271 sky130_fd_sc_hd__conb_1
X_13068_ clknet_leaf_167_clk _00535_ net1156 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08858__B total_design.core.ctrl.instruction\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12019_ total_design.lcd_display.row_2\[121\] _05848_ _05853_ total_design.lcd_display.row_2\[113\]
+ _05874_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12086__B1 _05812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07560_ total_design.core.regFile.register\[5\]\[19\] net807 net768 total_design.core.regFile.register\[7\]\[19\]
+ _03077_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__a221o_1
XANTENNA__08874__A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06511_ net742 net734 net730 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__and3_4
XANTENNA__08805__A1_N _02263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07491_ total_design.core.regFile.register\[20\]\[18\] net670 net604 total_design.core.regFile.register\[15\]\[18\]
+ _02998_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__a221o_1
XANTENNA__06665__Y _02233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11504__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09230_ net262 net2760 net456 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__mux2_1
X_06442_ _02013_ total_design.core.ctrl.instruction\[3\] _02012_ vssd1 vssd1 vccd1
+ vccd1 _02017_ sky130_fd_sc_hd__or3b_1
XFILLER_0_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ _04295_ _04299_ net330 vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06373_ total_design.core.ctrl.instruction\[24\] net918 _01948_ vssd1 vssd1 vccd1
+ vccd1 _01949_ sky130_fd_sc_hd__and3_1
XFILLER_0_161_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08112_ total_design.core.regFile.register\[20\]\[31\] net816 net814 total_design.core.regFile.register\[4\]\[31\]
+ net692 vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__a221o_1
XANTENNA__09909__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09092_ net314 _04337_ _04342_ net295 vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07804__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08043_ total_design.core.regFile.register\[23\]\[29\] net678 net612 total_design.core.regFile.register\[11\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold900 total_design.core.regFile.register\[15\]\[22\] vssd1 vssd1 vccd1 vccd1 net2216
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 total_design.core.regFile.register\[15\]\[18\] vssd1 vssd1 vccd1 vccd1 net2227
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 total_design.core.regFile.register\[2\]\[18\] vssd1 vssd1 vccd1 vccd1 net2238
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold933 total_design.core.regFile.register\[30\]\[10\] vssd1 vssd1 vccd1 vccd1 net2249
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 total_design.core.regFile.register\[27\]\[8\] vssd1 vssd1 vccd1 vccd1 net2260
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13728__Q total_design.core.data_bus_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold955 total_design.core.regFile.register\[9\]\[18\] vssd1 vssd1 vccd1 vccd1 net2271
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 total_design.core.regFile.register\[17\]\[27\] vssd1 vssd1 vccd1 vccd1 net2282
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold977 total_design.core.regFile.register\[7\]\[4\] vssd1 vssd1 vccd1 vccd1 net2293
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold988 total_design.core.regFile.register\[13\]\[31\] vssd1 vssd1 vccd1 vccd1 net2304
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ net261 net2378 net417 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__mux2_1
Xhold999 total_design.core.regFile.register\[16\]\[18\] vssd1 vssd1 vccd1 vccd1 net2315
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1118_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06240__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ _04185_ _04197_ _04198_ _04124_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout480_A _05011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06791__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08768__B _03595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ net337 _02868_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10810__C _05064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07827_ total_design.core.regFile.register\[18\]\[25\] net859 net836 total_design.core.regFile.register\[10\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout366_X net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07758_ total_design.core.regFile.register\[14\]\[23\] net624 net585 total_design.core.regFile.register\[28\]\[23\]
+ _03264_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__a221o_1
XANTENNA__08784__A _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06709_ total_design.core.regFile.register\[23\]\[3\] net679 net656 total_design.core.regFile.register\[29\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09493__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ total_design.core.regFile.register\[26\]\[22\] net870 net780 total_design.core.regFile.register\[27\]\[22\]
+ _03198_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09428_ net968 _02991_ net537 _02990_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09359_ _04505_ _04598_ net327 vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__mux2_1
XANTENNA__08048__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09819__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12370_ total_design.core.math.pc_val\[25\] net988 vssd1 vssd1 vccd1 vccd1 _01632_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11321_ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14040_ clknet_leaf_110_clk _01220_ net1225 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07008__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ _05399_ _05407_ _05500_ _05498_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__a31o_1
XANTENNA__12001__B1 _05838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10203_ _04542_ net2201 net390 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__mux2_1
X_11183_ _05441_ _05436_ _05434_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_128_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10134_ net230 net1965 net398 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10065_ net242 net2208 net406 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__mux2_1
XANTENNA__07192__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output128_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13824_ clknet_leaf_47_clk _01032_ net1097 vssd1 vssd1 vccd1 vccd1 total_design.core.data_access
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12068__B1 _05829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10967_ _05217_ _05225_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__nand2_1
XANTENNA__09484__A1 total_design.core.ctrl.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_97_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13755_ clknet_leaf_113_clk total_design.core.data_mem.stored_write_data\[30\] net1207
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12706_ clknet_leaf_129_clk _00173_ net1197 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13686_ clknet_leaf_50_clk total_design.core.data_mem.data_read_adr_i\[26\] net1099
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[26\] sky130_fd_sc_hd__dfrtp_1
X_10898_ _05151_ _05152_ _05153_ _05155_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__o22ai_4
XANTENNA__08039__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12637_ clknet_leaf_14_clk _00104_ net1026 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07247__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12568_ net1443 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06942__A total_design.core.ctrl.instruction\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_124_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11519_ net1726 _05630_ net152 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14307_ clknet_leaf_104_clk _00007_ net1238 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12499_ net979 total_design.core.instr_mem.instruction_i\[13\] vssd1 vssd1 vccd1
+ vccd1 _01704_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_117_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold207 total_design.lcd_display.row_1\[115\] vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold218 total_design.lcd_display.row_1\[111\] vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 total_design.lcd_display.row_1\[23\] vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ clknet_leaf_57_clk _01418_ net1119 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_169_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06380__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08747__B1 _02968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14169_ clknet_leaf_34_clk _01349_ net1068 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout709 net710 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08869__A _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09464__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06991_ net757 _02540_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[8\]
+ sky130_fd_sc_hd__and2_1
X_08730_ net944 net540 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.next_read
+ sky130_fd_sc_hd__or2_1
XANTENNA__10403__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11726__C net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08661_ total_design.lcd_display.cnt_500hz\[10\] _03941_ _03942_ vssd1 vssd1 vccd1
+ vccd1 _00006_ sky130_fd_sc_hd__o21a_1
XANTENNA__06525__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07612_ total_design.core.regFile.register\[3\]\[20\] net865 net758 total_design.core.regFile.register\[4\]\[20\]
+ _03125_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__a221o_1
X_08592_ _03904_ net880 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[13\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07543_ total_design.core.regFile.register\[5\]\[19\] net629 net605 total_design.core.regFile.register\[15\]\[19\]
+ _03045_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout159_A _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07486__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07474_ _02994_ _02995_ net721 vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06555__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09213_ net460 _04458_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__nand2_1
X_06425_ total_design.core.regFile.register\[10\]\[0\] net834 _01975_ _01944_ _01955_
+ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_134_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09144_ _01746_ _02391_ _02392_ _04101_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07238__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06356_ _01928_ _01931_ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__nor2_8
XFILLER_0_133_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09075_ _04324_ _04325_ net329 vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__mux2_1
X_06287_ net930 _01863_ _01865_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1235_A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08026_ total_design.core.regFile.register\[28\]\[29\] net853 net802 total_design.core.regFile.register\[8\]\[29\]
+ _03521_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold730 total_design.core.regFile.register\[5\]\[27\] vssd1 vssd1 vccd1 vccd1 net2046
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 total_design.core.regFile.register\[17\]\[3\] vssd1 vssd1 vccd1 vccd1 net2057
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 total_design.core.regFile.register\[2\]\[6\] vssd1 vssd1 vccd1 vccd1 net2068
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 total_design.core.regFile.register\[3\]\[2\] vssd1 vssd1 vccd1 vccd1 net2079
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 total_design.core.regFile.register\[2\]\[29\] vssd1 vssd1 vccd1 vccd1 net2090
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold785 total_design.core.regFile.register\[29\]\[0\] vssd1 vssd1 vccd1 vccd1 net2101
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 total_design.core.regFile.register\[5\]\[19\] vssd1 vssd1 vccd1 vccd1 net2112
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09977_ net187 net2273 net419 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout862_A net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06764__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10313__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ _04180_ _04181_ net459 vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1430 total_design.core.regFile.register\[18\]\[6\] vssd1 vssd1 vccd1 vccd1 net2746
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 total_design.core.regFile.register\[30\]\[9\] vssd1 vssd1 vccd1 vccd1 net2757
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14289__Q net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1452 total_design.core.regFile.register\[9\]\[6\] vssd1 vssd1 vccd1 vccd1 net2768
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1463 total_design.core.regFile.register\[19\]\[17\] vssd1 vssd1 vccd1 vccd1 net2779
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08859_ total_design.core.ctrl.instruction\[9\] total_design.core.ctrl.instruction\[10\]
+ net556 vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__nand3_2
Xhold1474 total_design.core.regFile.register\[10\]\[7\] vssd1 vssd1 vccd1 vccd1 net2790
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1485 total_design.core.regFile.register\[14\]\[22\] vssd1 vssd1 vccd1 vccd1 net2801
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11870_ _05752_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__inv_2
Xhold1496 total_design.core.regFile.register\[19\]\[30\] vssd1 vssd1 vccd1 vccd1 net2812
+ sky130_fd_sc_hd__dlygate4sd3_1
X_10821_ _05063_ _05074_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07477__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10752_ net2869 net355 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__and2_1
X_13540_ clknet_leaf_107_clk _01007_ net1223 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[0\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14248__RESET_B net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13471_ clknet_leaf_183_clk _00938_ net1040 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14550__1270 vssd1 vssd1 vccd1 vccd1 _14550__1270/HI net1270 sky130_fd_sc_hd__conb_1
X_10683_ net190 net2330 net362 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12422_ net900 _03602_ net524 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__a21o_1
XANTENNA__07229__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12353_ _01613_ _01614_ _01616_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__or3_1
XANTENNA__06481__B net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11304_ _05514_ _05520_ _05554_ _05558_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12284_ total_design.core.math.pc_val\[16\] total_design.core.program_count.imm_val_reg\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_75_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14023_ clknet_leaf_82_clk _01203_ net1241 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11235_ _05490_ _05493_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_147_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07401__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ net514 _05184_ _05424_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10731__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06755__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ net167 net2812 net404 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__mux2_1
XANTENNA__12289__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10223__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11097_ net513 _05220_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__and2_2
XFILLER_0_101_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10048_ net172 net2515 net411 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_160_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold90 total_design.keypad0.counter\[18\] vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06937__A _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07180__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13807_ clknet_leaf_71_clk total_design.core.data_mem.data_cpu_i\[16\] net1211 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[16\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09457__A1 _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11999_ total_design.lcd_display.row_2\[96\] _05846_ _05850_ total_design.lcd_display.row_2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_11_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09032__B _04283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13738_ clknet_leaf_77_clk total_design.core.data_mem.stored_write_data\[13\] net1214
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_128_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06375__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13669_ clknet_leaf_63_clk total_design.core.data_mem.data_read_adr_i\[9\] net1125
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06210_ _01788_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07190_ total_design.core.regFile.register\[30\]\[12\] net840 net806 total_design.core.regFile.register\[5\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a22o_1
XANTENNA__06672__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06141_ total_design.lcd_display.currentState\[0\] vssd1 vssd1 vccd1 vccd1 _01724_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07640__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09900_ net221 net2555 net427 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__mux2_1
XANTENNA__10527__A0 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout506 net507 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__buf_4
XFILLER_0_1_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09393__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout517 net519 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__clkbuf_4
X_09831_ net225 total_design.core.regFile.register\[27\]\[15\] net437 vssd1 vssd1
+ vccd1 vccd1 _00150_ sky130_fd_sc_hd__mux2_1
Xfanout528 _06017_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_2
Xfanout539 _03676_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10133__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09762_ net235 net2151 net443 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__mux2_1
X_06974_ total_design.core.regFile.register\[24\]\[8\] net792 net788 total_design.core.regFile.register\[13\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__a22o_1
XANTENNA__09922__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08713_ total_design.keypad0.counter\[3\] total_design.keypad0.counter\[4\] _03950_
+ total_design.keypad0.counter\[5\] vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__a31o_1
X_09693_ net472 _03506_ _04264_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout276_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ total_design.lcd_display.cnt_500hz\[3\] _03921_ total_design.lcd_display.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07171__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08575_ net1839 net338 net718 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[30\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__13741__Q total_design.core.data_bus_o\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout443_A _04969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1185_A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07526_ _03038_ _03039_ _03036_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__a21boi_4
XANTENNA__07459__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07457_ total_design.core.regFile.register\[22\]\[17\] net775 net758 total_design.core.regFile.register\[4\]\[17\]
+ _02975_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout610_A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08781__B _02770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06408_ net923 net947 net909 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07388_ total_design.core.regFile.register\[19\]\[16\] net642 net568 total_design.core.regFile.register\[12\]\[16\]
+ _02898_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09127_ _02341_ _04350_ _04375_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__a21oi_1
X_06339_ total_design.core.ctrl.instruction\[2\] total_design.core.ctrl.instruction\[3\]
+ total_design.core.ctrl.instruction\[0\] total_design.core.ctrl.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__or4bb_4
XANTENNA__09620__A1 _03421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10308__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10766__B1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07631__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09058_ net322 _04307_ _04309_ net312 vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__a211o_1
XFILLER_0_103_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11487__X _05682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__A2 total_design.core.data_mem.data_cpu_i\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08009_ total_design.core.regFile.register\[0\]\[28\] net684 _03502_ _03505_ vssd1
+ vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_92_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10781__A3 total_design.core.data_bus_o\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold560 total_design.core.mem_ctrl.state\[1\] vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold571 total_design.keypad0.key_counter\[0\] vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ net350 _05278_ _05268_ _05266_ _05264_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_124_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold582 total_design.core.regFile.register\[29\]\[30\] vssd1 vssd1 vccd1 vccd1 net1898
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 total_design.core.regFile.register\[26\]\[2\] vssd1 vssd1 vccd1 vccd1 net1909
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06737__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_X net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13223__RESET_B net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10043__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09832__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ clknet_leaf_107_clk _00438_ net1224 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1260 total_design.core.regFile.register\[9\]\[24\] vssd1 vssd1 vccd1 vccd1 net2576
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 total_design.core.regFile.register\[20\]\[7\] vssd1 vssd1 vccd1 vccd1 net2587
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ _05796_ total_design.keypad0.key_out\[3\] net530 vssd1 vssd1 vccd1 vccd1
+ _01450_ sky130_fd_sc_hd__mux2_1
XANTENNA__11494__A1 _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1282 total_design.core.regFile.register\[17\]\[18\] vssd1 vssd1 vccd1 vccd1 net2598
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1293 total_design.core.regFile.register\[22\]\[16\] vssd1 vssd1 vccd1 vccd1 net2609
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07162__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11853_ _05727_ _05728_ _05738_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_68_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06476__B net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10804_ net521 _05062_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__nand2_2
X_11784_ net929 _01810_ _05694_ net953 net1506 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__a32o_1
XFILLER_0_138_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13523_ clknet_leaf_179_clk _00990_ net1041 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10735_ total_design.core.regFile.register\[0\]\[10\] net353 vssd1 vssd1 vccd1 vccd1
+ _01009_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11602__S net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13454_ clknet_leaf_190_clk _00921_ net1034 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10666_ net265 net1948 net361 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__mux2_1
XANTENNA__10726__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14482__Q total_design.core.ctrl.instruction\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_201_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12405_ net900 _03512_ net525 vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10218__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13385_ clknet_leaf_18_clk _00852_ net1046 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10597_ net282 net2733 net365 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10221__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__clkbuf_4
X_12336_ net990 _01599_ _01600_ _01601_ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06976__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12267_ _06098_ _06099_ _06100_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12433__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11218_ _05471_ _05476_ _05355_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a21o_2
X_14006_ clknet_leaf_111_clk _01186_ net1210 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12198_ _06037_ _06046_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__nand2_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_162_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_128_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11149_ _05399_ _05407_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11485__A1 _05651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07770__B _03273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07689__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06690_ total_design.core.regFile.register\[4\]\[3\] net815 _02254_ _02255_ _02256_
+ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06667__A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06900__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08360_ _03713_ _03716_ _03718_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__and3_2
XFILLER_0_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07311_ _02791_ _02841_ _02842_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__or3_1
XANTENNA__11788__A2 _01847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08291_ total_design.core.data_mem.data_write_adr_reg\[3\] net549 net541 total_design.core.data_mem.data_read_adr_reg\[3\]
+ net945 vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06673__Y _02241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11512__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07242_ total_design.core.regFile.register\[25\]\[13\] net845 net770 total_design.core.regFile.register\[7\]\[13\]
+ _02777_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07173_ total_design.core.regFile.register\[29\]\[12\] net655 net633 total_design.core.regFile.register\[16\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__a22o_1
XANTENNA__10128__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06552__D net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13734__RESET_B net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07613__B1 _01992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06967__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09366__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout303 _05458_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_4
XANTENNA__09218__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout314 net315 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_2
XANTENNA__13736__Q total_design.core.data_bus_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout325 net327 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_1
XANTENNA__06719__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 net337 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_2
Xfanout347 _01685_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__buf_4
X_09814_ total_design.core.ctrl.instruction\[7\] total_design.core.ctrl.instruction\[8\]
+ net556 vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__nand3_2
Xfanout358 _05017_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_4
Xfanout369 _05013_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_8
XANTENNA__09118__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07392__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__X _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ net161 net2356 net455 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout560_A _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09669__A1 _03512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06957_ total_design.core.regFile.register\[19\]\[8\] net642 _02505_ _02506_ _02507_
+ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11476__A1 _05609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06888_ net721 _02398_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__nor2_1
X_09676_ _04687_ _04731_ _04897_ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__o211a_1
XANTENNA__07144__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08627_ total_design.lcd_display.cnt_500hz\[1\] total_design.lcd_display.cnt_500hz\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout825_A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ net717 _03904_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[13\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07509_ total_design.core.regFile.register\[19\]\[18\] net823 net783 total_design.core.regFile.register\[2\]\[18\]
+ _03018_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__a221o_1
X_08489_ total_design.data_in_BUS\[7\] _01888_ _03841_ net519 vssd1 vssd1 vccd1 vccd1
+ _03842_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout613_X net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11422__S net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10520_ net182 net2470 net482 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07852__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ net194 net2120 net381 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10038__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08016__B _03512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13170_ clknet_leaf_145_clk _00637_ net1179 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07604__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09827__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10382_ net205 net2513 net484 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout982_X net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12121_ total_design.lcd_display.row_1\[70\] _05804_ _05849_ total_design.lcd_display.row_2\[54\]
+ _05971_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__a221o_1
XANTENNA__06958__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13404__RESET_B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12052_ total_design.lcd_display.currentState\[3\] _05751_ net474 _05746_ vssd1 vssd1
+ vccd1 vccd1 _05911_ sky130_fd_sc_hd__o211a_1
Xhold390 total_design.lcd_display.row_2\[6\] vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ _05244_ _05245_ _05256_ _05261_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07383__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 net872 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__clkbuf_8
Xfanout881 net882 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__clkbuf_4
Xfanout892 net893 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11467__A1 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10501__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ clknet_leaf_132_clk _00421_ net1200 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1090 net111 vssd1 vssd1 vccd1 vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07135__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_107_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14477__Q total_design.core.ctrl.instruction\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _05781_ _05782_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_29_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_193_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_193_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12885_ clknet_leaf_167_clk _00352_ net1155 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11836_ total_design.lcd_display.currentState\[0\] _05719_ vssd1 vssd1 vccd1 vccd1
+ _05723_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14555_ net1275 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XANTENNA__08096__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ net930 _01904_ _05697_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_155_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_140_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13506_ clknet_leaf_130_clk _00973_ net1198 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10718_ net181 net2542 net359 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__mux2_1
X_14486_ clknet_leaf_32_clk _01553_ net1063 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_130_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11698_ net33 net935 net878 net1679 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13437_ clknet_leaf_11_clk _00904_ net1025 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10649_ net194 net2423 net476 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13368_ clknet_leaf_138_clk _00835_ net1185 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_155_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06949__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ net899 _03090_ net522 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13299_ clknet_leaf_179_clk _00766_ net1034 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07860_ total_design.core.regFile.register\[14\]\[25\] net625 net578 total_design.core.regFile.register\[27\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__a22o_1
XANTENNA__08020__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07374__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06811_ total_design.core.regFile.register\[17\]\[5\] net821 _02369_ _02370_ vssd1
+ vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07791_ total_design.core.regFile.register\[16\]\[24\] net855 net765 total_design.core.regFile.register\[6\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11507__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11458__A1 _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09530_ _04744_ _04761_ _03230_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__o21a_1
X_06742_ total_design.core.regFile.register\[26\]\[4\] net869 net767 total_design.core.regFile.register\[7\]\[4\]
+ _02293_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10411__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07126__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ total_design.core.ctrl.instruction\[18\] net886 net754 total_design.core.data_cpu_o\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__a22o_1
X_06673_ _02213_ _02240_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__xnor2_4
Xclkbuf_leaf_184_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_184_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08412_ _03767_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09392_ _04194_ _04624_ _04626_ _04159_ _04628_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08343_ total_design.core.data_mem.data_write_adr_reg\[29\] net547 net539 total_design.core.data_mem.data_read_adr_reg\[29\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08087__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout141_A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08274_ net1484 net558 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[24\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_15_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07834__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07225_ total_design.core.regFile.register\[30\]\[13\] net659 net640 total_design.core.regFile.register\[19\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout406_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1050_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07156_ total_design.core.ctrl.instruction\[12\] _02641_ vssd1 vssd1 vccd1 vccd1
+ _02696_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10197__A1 _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07087_ total_design.core.regFile.register\[0\]\[10\] net873 _02625_ _02631_ vssd1
+ vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_140_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09339__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1109 net1121 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout775_A _01990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout133 _05686_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_4
Xfanout144 _05684_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_2
Xfanout155 _05681_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_4
Xfanout166 _04950_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_35_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout177 net179 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__buf_1
Xfanout188 _04843_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout942_A _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_2
X_07989_ _03486_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i\[28\]
+ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout563_X net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11449__A1 _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10321__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09728_ _03596_ _03597_ _04933_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07117__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12110__A2 _05804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ total_design.core.math.pc_val\[27\] _04861_ vssd1 vssd1 vccd1 vccd1 _04886_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_26_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_175_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_175_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08865__A2 total_design.core.ctrl.instruction\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12670_ clknet_leaf_181_clk _00137_ net1044 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11621_ _05621_ net1851 net133 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__mux2_1
XANTENNA__08078__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14340_ clknet_leaf_67_clk _01501_ net1112 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_13_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11552_ net1567 _05630_ net147 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06473__C net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10503_ net249 net2320 net483 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__mux2_1
X_11483_ net1555 _05633_ net154 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14271_ net986 _01447_ net1085 vssd1 vssd1 vccd1 vccd1 total_design.data_from_keypad\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09027__C1 _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13222_ clknet_leaf_194_clk _00689_ net1011 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10434_ net273 net2768 net383 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10365_ net268 net2536 net486 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__mux2_1
X_13153_ clknet_leaf_126_clk _00620_ net1192 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ total_design.lcd_display.row_2\[29\] _05832_ net348 total_design.lcd_display.row_2\[61\]
+ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__a22o_1
X_13084_ clknet_leaf_29_clk _00551_ net1073 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10296_ net285 net2374 net492 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__mux2_1
X_12035_ total_design.lcd_display.row_1\[66\] _05804_ _05821_ total_design.lcd_display.row_1\[42\]
+ _05892_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08002__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09750__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07356__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07761__C1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10231__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09305__B net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13986_ clknet_leaf_85_clk _01166_ net1247 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07108__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12101__A2 _05814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12937_ clknet_leaf_17_clk _00404_ net1046 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_166_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_166_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_157_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ clknet_leaf_105_clk _00335_ net1233 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08069__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11819_ _05711_ net1859 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_174_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ clknet_leaf_183_clk _00266_ net1039 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14538_ net1310 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_0_141_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06383__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14469_ clknet_leaf_54_clk net1389 net1110 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07010_ total_design.core.regFile.register\[18\]\[9\] net610 net568 total_design.core.regFile.register\[12\]\[9\]
+ _02557_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10406__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07595__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08961_ net462 _04212_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07912_ total_design.core.regFile.register\[11\]\[26\] net613 _03407_ _03410_ _03412_
+ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__a2111o_1
X_08892_ net469 _02334_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__nor2_1
XANTENNA__07347__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ total_design.core.regFile.register\[13\]\[25\] net787 _03331_ _03346_ vssd1
+ vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10141__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ _03254_ _03279_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__or2_2
XFILLER_0_116_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09930__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09513_ _03187_ net705 _04745_ net536 vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__a211oi_1
XANTENNA__06558__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06725_ _02286_ net314 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_157_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_157_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout356_A _05018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06656_ total_design.core.regFile.register\[26\]\[2\] net644 net612 total_design.core.regFile.register\[11\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__a22o_1
X_09444_ net506 _04680_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_82_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_166_Right_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09231__A _02515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06587_ total_design.core.regFile.register\[2\]\[1\] net740 net737 net731 vssd1 vssd1
+ vccd1 vccd1 _02158_ sky130_fd_sc_hd__and4_1
X_09375_ net506 _04614_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout144_X net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1265_A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08326_ net1477 net938 _03697_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[20\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07807__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08257_ net1365 net559 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[7\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_117_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07208_ _02742_ _02745_ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__xnor2_4
Xclkbuf_3_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08188_ net891 _03646_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[31\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07139_ total_design.core.regFile.register\[25\]\[11\] net842 net789 total_design.core.regFile.register\[13\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__a22o_1
XANTENNA__10316__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07586__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ net171 net2694 net398 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06794__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ net177 net2033 net407 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07743__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06749__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ clknet_leaf_58_clk _01048_ net1119 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_stored\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10051__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09840__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__Y _05804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13771_ clknet_leaf_58_clk total_design.core.data_mem.stored_data_adr\[14\] net1118
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[14\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_148_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_148_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10983_ _05241_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12722_ clknet_leaf_139_clk _00189_ net1184 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07510__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11390__B _05645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ clknet_leaf_7_clk _00120_ net1016 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06484__B net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11604_ _05657_ net1717 net138 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12584_ clknet_leaf_171_clk _00051_ net1056 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14323_ clknet_leaf_68_clk _01484_ net1111 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_52_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11535_ net1660 _05655_ net145 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11610__S net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14254_ clknet_leaf_104_clk _01434_ net1234 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11466_ net1615 _05670_ net155 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10734__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14490__Q total_design.core.ctrl.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13205_ clknet_leaf_158_clk _00672_ net1141 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10417_ net197 net1994 net386 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14185_ clknet_leaf_79_clk _01365_ net1218 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
X_11397_ total_design.core.data_bus_o\[17\] net699 _05573_ vssd1 vssd1 vccd1 vccd1
+ _05656_ sky130_fd_sc_hd__a21oi_2
X_13136_ clknet_leaf_186_clk _00603_ net1031 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10348_ net210 net2180 net489 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__mux2_1
XANTENNA__11846__A _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12441__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10279_ net221 net2453 net499 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__mux2_1
X_13067_ clknet_leaf_107_clk _00534_ net1224 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07329__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12018_ total_design.lcd_display.row_2\[73\] _05806_ _05830_ total_design.lcd_display.row_1\[1\]
+ _05878_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__a221o_1
XANTENNA__06537__A0 total_design.core.data_mem.data_cpu_i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09750__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06378__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13969_ clknet_leaf_95_clk _01149_ net1256 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[51\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_139_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_139_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06510_ total_design.core.regFile.register\[28\]\[0\] net747 net739 net727 vssd1
+ vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__and4_1
XANTENNA__08874__B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07490_ total_design.core.regFile.register\[8\]\[18\] net593 net589 total_design.core.regFile.register\[1\]\[18\]
+ _03000_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_17_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07501__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08593__C net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06441_ _02013_ _01735_ _02012_ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__and3b_2
XFILLER_0_75_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09160_ net323 _04293_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06372_ net951 net950 net966 net965 net952 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_174_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11597__A0 _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08111_ total_design.core.regFile.register\[16\]\[31\] net855 net847 total_design.core.regFile.register\[15\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09091_ net328 _04339_ _04340_ _04341_ net318 vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08042_ total_design.core.regFile.register\[29\]\[29\] net655 net589 total_design.core.regFile.register\[1\]\[29\]
+ _03534_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__a221o_1
Xhold901 total_design.data_in_BUS\[16\] vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 total_design.core.regFile.register\[10\]\[15\] vssd1 vssd1 vccd1 vccd1 net2228
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold923 total_design.core.regFile.register\[6\]\[1\] vssd1 vssd1 vccd1 vccd1 net2239
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 total_design.core.regFile.register\[1\]\[19\] vssd1 vssd1 vccd1 vccd1 net2250
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10136__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold945 total_design.core.regFile.register\[15\]\[2\] vssd1 vssd1 vccd1 vccd1 net2261
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold956 total_design.core.regFile.register\[24\]\[24\] vssd1 vssd1 vccd1 vccd1 net2272
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09925__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08765__A1 _03395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold967 total_design.core.regFile.register\[20\]\[24\] vssd1 vssd1 vccd1 vccd1 net2283
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 total_design.core.regFile.register\[2\]\[3\] vssd1 vssd1 vccd1 vccd1 net2294
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 total_design.keypad0.key_counter\[1\] vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ net267 net2727 net415 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06240__A2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08944_ _04158_ _04184_ _04191_ _04157_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ net470 _02818_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_32_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout473_A _02111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07826_ net749 _03330_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[24\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07017__Y _02565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07740__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ total_design.core.regFile.register\[10\]\[23\] net616 net577 total_design.core.regFile.register\[27\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout640_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08784__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06708_ total_design.core.regFile.register\[25\]\[3\] net648 net571 total_design.core.regFile.register\[17\]\[3\]
+ _02271_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07688_ total_design.core.regFile.register\[24\]\[22\] net791 net768 total_design.core.regFile.register\[7\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13248__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ net313 _02337_ _04104_ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__or3_4
X_06639_ _02191_ _02192_ _02207_ _02208_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__or4_1
XFILLER_0_109_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09358_ _04597_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__inv_2
XANTENNA__09245__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08309_ total_design.core.data_mem.data_write_adr_reg\[12\] net548 net540 total_design.core.data_mem.data_read_adr_reg\[12\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10835__A total_design.core.data_bus_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09289_ net315 _04326_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11430__S net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11320_ _05494_ _05495_ _05481_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_16_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout895_X net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11251_ _05500_ _05506_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10046__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10012__A0 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07559__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10202_ net256 net2599 net389 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__mux2_1
XANTENNA__09835__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11182_ _05431_ _05436_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10133_ net236 net2556 net399 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input34_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10064_ net254 net2818 net406 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__mux2_1
XANTENNA__06479__B net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07192__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823_ clknet_leaf_44_clk _01031_ net1087 vssd1 vssd1 vccd1 vccd1 total_design.core.mem_ctrl.next_next_fetch
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09469__C1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11605__S net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13671__RESET_B net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13754_ clknet_leaf_113_clk total_design.core.data_mem.stored_write_data\[29\] net1207
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[29\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_168_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10966_ _05221_ _05222_ _05218_ _05219_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10729__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12705_ clknet_leaf_121_clk _00172_ net1167 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06298__A2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13685_ clknet_leaf_51_clk total_design.core.data_mem.data_read_adr_i\[25\] net1093
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10897_ _05153_ _05155_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12636_ clknet_leaf_30_clk _00103_ net1060 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11579__A0 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09236__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12567_ net1425 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12436__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07798__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14306_ clknet_leaf_104_clk _00006_ net1236 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11518_ net1835 _05651_ net149 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12498_ net977 total_design.core.ctrl.instruction\[12\] net882 _01703_ vssd1 vssd1
+ vccd1 vccd1 _01551_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_117_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold208 total_design.lcd_display.row_1\[108\] vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold219 total_design.lcd_display.row_1\[69\] vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14237_ clknet_leaf_57_clk _01417_ net1119 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11449_ net1575 _05646_ net158 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09745__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08747__B2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14168_ clknet_leaf_34_clk _01348_ net1066 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06758__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13119_ clknet_leaf_183_clk _00586_ net1040 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_84_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14099_ clknet_leaf_93_clk _01279_ net1257 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[53\]
+ sky130_fd_sc_hd__dfrtp_1
X_06990_ _02496_ _02539_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__xor2_2
XANTENNA__07970__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09172__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ total_design.lcd_display.cnt_500hz\[10\] _03941_ net711 vssd1 vssd1 vccd1
+ vccd1 _03942_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_79_1092 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07183__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07611_ total_design.core.regFile.register\[12\]\[20\] _01980_ net782 total_design.core.regFile.register\[27\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__a22o_1
X_08591_ _03901_ net880 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[12\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06930__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11515__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07542_ total_design.core.regFile.register\[30\]\[19\] net660 net594 total_design.core.regFile.register\[8\]\[19\]
+ _03059_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_93_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07473_ total_design.core.ctrl.instruction\[18\] _02945_ vssd1 vssd1 vccd1 vccd1
+ _02995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09212_ net469 _02515_ _04144_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__o21a_1
XANTENNA__06555__D net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06424_ total_design.core.regFile.register\[21\]\[0\] net928 net910 net908 vssd1
+ vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__and4_1
XFILLER_0_174_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09143_ _02391_ _04188_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__nand2_1
X_06355_ net951 net950 _01930_ net952 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__o211a_2
XANTENNA__07789__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ _04251_ _04255_ net468 vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__mux2_1
X_06286_ total_design.core.data_adr_o\[7\] _01864_ net964 vssd1 vssd1 vccd1 vccd1
+ _01865_ sky130_fd_sc_hd__mux2_1
XANTENNA__13739__Q total_design.core.data_bus_o\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06997__B1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08025_ total_design.core.regFile.register\[3\]\[29\] net865 net831 total_design.core.regFile.register\[31\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1130_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold720 total_design.core.regFile.register\[19\]\[25\] vssd1 vssd1 vccd1 vccd1 net2036
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 total_design.core.regFile.register\[5\]\[5\] vssd1 vssd1 vccd1 vccd1 net2047
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 total_design.core.regFile.register\[23\]\[6\] vssd1 vssd1 vccd1 vccd1 net2058
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1228_A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold753 total_design.core.regFile.register\[9\]\[15\] vssd1 vssd1 vccd1 vccd1 net2069
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12534__A2 total_design.core.ctrl.instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold764 total_design.core.regFile.register\[11\]\[5\] vssd1 vssd1 vccd1 vccd1 net2080
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 total_design.core.regFile.register\[26\]\[18\] vssd1 vssd1 vccd1 vccd1 net2091
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 total_design.core.regFile.register\[11\]\[4\] vssd1 vssd1 vccd1 vccd1 net2102
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08779__B total_design.core.data_mem.data_cpu_i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold797 total_design.core.regFile.register\[17\]\[23\] vssd1 vssd1 vccd1 vccd1 net2113
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ net190 net2246 net419 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07961__A2 total_design.core.data_mem.data_cpu_i\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08927_ _02917_ _02968_ net470 vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout855_A _01947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1420 total_design.core.regFile.register\[18\]\[9\] vssd1 vssd1 vccd1 vccd1 net2736
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1431 total_design.core.regFile.register\[20\]\[17\] vssd1 vssd1 vccd1 vccd1 net2747
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1442 total_design.core.regFile.register\[22\]\[26\] vssd1 vssd1 vccd1 vccd1 net2758
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08858_ total_design.core.ctrl.instruction\[7\] total_design.core.ctrl.instruction\[8\]
+ _04111_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__nand3b_2
XANTENNA__07174__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1453 total_design.core.regFile.register\[10\]\[9\] vssd1 vssd1 vccd1 vccd1 net2769
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 total_design.core.regFile.register\[3\]\[8\] vssd1 vssd1 vccd1 vccd1 net2780
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1475 total_design.core.regFile.register\[5\]\[31\] vssd1 vssd1 vccd1 vccd1 net2791
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1486 total_design.core.regFile.register\[19\]\[24\] vssd1 vssd1 vccd1 vccd1 net2802
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07809_ total_design.core.regFile.register\[13\]\[24\] net667 _03311_ _03312_ _03313_
+ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__a2111o_1
Xhold1497 total_design.core.regFile.register\[3\]\[20\] vssd1 vssd1 vccd1 vccd1 net2813
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06921__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08789_ _02868_ total_design.core.data_mem.data_cpu_i\[15\] vssd1 vssd1 vccd1 vccd1
+ _04044_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_140_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11425__S net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10820_ net521 _05078_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10751_ total_design.core.regFile.register\[0\]\[26\] net355 vssd1 vssd1 vccd1 vccd1
+ _01025_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_49_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout810_X net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13470_ clknet_leaf_157_clk _00937_ net1141 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10682_ net196 net2392 net361 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12421_ net993 _04946_ _01677_ net895 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12352_ total_design.core.math.pc_val\[23\] net988 vssd1 vssd1 vccd1 vccd1 _01616_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10784__A1 total_design.core.data_bus_o\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11303_ _05560_ _05561_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_75_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12283_ total_design.core.math.pc_val\[16\] total_design.core.program_count.imm_val_reg\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14022_ clknet_leaf_100_clk _01202_ net1236 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_11234_ _05391_ _05395_ _05397_ _05489_ _05491_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_147_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11165_ _05411_ _05418_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10504__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07952__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10116_ net170 net2020 net402 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__mux2_1
X_11096_ net513 _05291_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__nand2_1
X_10047_ net177 net2531 net411 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07165__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 total_design.core.data_mem.data_cpu_i_reg\[16\] vssd1 vssd1 vccd1 vccd1 net1396
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_160_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold91 total_design.core.data_mem.data_bus_i_reg\[26\] vssd1 vssd1 vccd1 vccd1 net1407
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07704__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06912__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13806_ clknet_leaf_71_clk total_design.core.data_mem.data_cpu_i\[15\] net1209 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[15\] sky130_fd_sc_hd__dfrtp_1
X_11998_ total_design.lcd_display.row_2\[40\] _05844_ _05849_ total_design.lcd_display.row_2\[48\]
+ _05854_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13737_ clknet_leaf_76_clk total_design.core.data_mem.stored_write_data\[12\] net1214
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[12\] sky130_fd_sc_hd__dfrtp_1
X_10949_ _05124_ _05207_ _05057_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13668_ clknet_leaf_66_clk total_design.core.data_mem.data_read_adr_i\[8\] net1122
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11016__A2 _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12619_ clknet_leaf_127_clk _00086_ net1191 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06691__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13599_ clknet_leaf_61_clk net1349 net1129 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06672__B net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10224__A0 _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06140_ total_design.lcd_display.currentState\[4\] vssd1 vssd1 vccd1 vccd1 _01723_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_27_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10194__B net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06979__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06391__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12516__A2 total_design.core.ctrl.instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ net234 net2820 net435 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__mux2_1
Xfanout507 _04122_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_8
Xfanout518 net519 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10414__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout529 _05787_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__buf_2
XANTENNA__07943__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09761_ net228 net2314 net443 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06973_ total_design.core.regFile.register\[30\]\[8\] net840 net766 total_design.core.regFile.register\[6\]\[8\]
+ _02523_ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__a221o_1
XANTENNA__09145__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08712_ _03953_ _03975_ _03976_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__nor3_1
X_09692_ _03557_ net509 net448 _03554_ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__o221a_1
XANTENNA__09504__A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ total_design.lcd_display.cnt_500hz\[3\] total_design.lcd_display.cnt_500hz\[4\]
+ _03921_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__and3_1
XANTENNA__06903__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08574_ total_design.data_in_BUS\[29\] net341 net719 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[29\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_166_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07525_ total_design.core.ctrl.instruction\[31\] net885 _02149_ _03043_ net550 vssd1
+ vssd1 vccd1 vccd1 total_design.core.ctrl.imm_32\[19\] sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1080_A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_61_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout436_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08120__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1178_A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07456_ _02976_ _02977_ _02978_ _02979_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_79_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06407_ total_design.core.regFile.register\[24\]\[0\] net928 net919 net915 vssd1
+ vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__and4_1
XFILLER_0_174_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06682__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07387_ total_design.core.regFile.register\[27\]\[16\] net579 _02913_ net688 vssd1
+ vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout603_A _02076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09126_ _02335_ _02338_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__nor2_1
X_06338_ total_design.core.ctrl.instruction\[2\] total_design.core.ctrl.instruction\[3\]
+ total_design.core.ctrl.instruction\[0\] total_design.core.ctrl.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_17_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06269_ total_design.core.instr_mem.instruction_adr_i\[10\] total_design.core.instr_mem.instruction_adr_stored\[10\]
+ net985 vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__mux2_1
X_09057_ net462 _04148_ _04308_ net324 vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1133_X net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08008_ _03489_ _03492_ _03494_ _03504_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_92_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold550 total_design.data_in_BUS\[8\] vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 total_design.core.regFile.register\[6\]\[0\] vssd1 vssd1 vccd1 vccd1 net1877
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout593_X net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold572 total_design.core.regFile.register\[24\]\[1\] vssd1 vssd1 vccd1 vccd1 net1888
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 total_design.core.regFile.register\[14\]\[6\] vssd1 vssd1 vccd1 vccd1 net1899
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10324__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 total_design.core.regFile.register\[30\]\[2\] vssd1 vssd1 vccd1 vccd1 net1910
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07934__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ net265 net2537 net421 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout858_X net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ clknet_leaf_22_clk _00437_ net1055 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[18\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07147__B1 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1250 total_design.core.regFile.register\[8\]\[23\] vssd1 vssd1 vccd1 vccd1 net2566
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 total_design.core.regFile.register\[19\]\[26\] vssd1 vssd1 vccd1 vccd1 net2577
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11921_ _03907_ _05779_ net38 vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a21o_1
Xhold1272 total_design.core.regFile.register\[22\]\[10\] vssd1 vssd1 vccd1 vccd1 net2588
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1283 total_design.core.regFile.register\[16\]\[10\] vssd1 vssd1 vccd1 vccd1 net2599
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1294 total_design.core.regFile.register\[30\]\[24\] vssd1 vssd1 vccd1 vccd1 net2610
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11852_ total_design.lcd_display.currentState\[1\] total_design.lcd_display.currentState\[2\]
+ total_design.lcd_display.currentState\[0\] vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06249__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ total_design.core.data_bus_o\[10\] net699 vssd1 vssd1 vccd1 vccd1 _05062_
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_138_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11950__Y _05812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11783_ net929 _01813_ _05694_ net953 net1508 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_52_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08972__B _02666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08111__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07869__A _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13522_ clknet_leaf_139_clk _00989_ net1183 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10734_ total_design.core.regFile.register\[0\]\[9\] net356 vssd1 vssd1 vccd1 vccd1
+ _01008_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06773__A _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13453_ clknet_leaf_6_clk _00920_ net1017 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10665_ net275 net2068 net363 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__mux2_1
XANTENNA__08036__Y _03532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_149_Left_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12404_ net991 _01660_ _01661_ _01662_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13384_ clknet_leaf_170_clk _00851_ net1159 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10596_ net268 total_design.core.regFile.register\[4\]\[3\] net366 vssd1 vssd1 vccd1
+ vccd1 _00874_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12335_ net990 _04756_ net894 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_11_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06425__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12266_ total_design.core.math.pc_val\[14\] total_design.core.program_count.imm_val_reg\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10742__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14005_ clknet_leaf_91_clk _01185_ net1262 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11217_ net302 _05473_ _05474_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__and3_1
XANTENNA__10234__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__clkbuf_4
X_12197_ total_design.core.math.pc_val\[4\] total_design.core.program_count.imm_val_reg\[4\]
+ total_design.core.program_count.imm_val_reg\[5\] total_design.core.math.pc_val\[5\]
+ _06030_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07386__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_162_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07925__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__clkbuf_4
X_11148_ _05402_ _05403_ _05405_ _05358_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_158_Left_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11079_ _05290_ _05292_ _05285_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__a21o_1
XANTENNA__07138__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12131__B1 _05829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09324__A _02718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10693__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06667__B total_design.core.ctrl.imm_32\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06386__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_43_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08882__B _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07310_ _02689_ _02743_ _02744_ _02793_ _02739_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__o311a_1
X_08290_ net1471 net940 _03679_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[2\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_167_Left_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07241_ total_design.core.regFile.register\[26\]\[13\] net869 net819 total_design.core.regFile.register\[17\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__a22o_1
XANTENNA__10409__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07172_ total_design.core.regFile.register\[2\]\[12\] net639 net623 total_design.core.regFile.register\[4\]\[12\]
+ _02710_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__a221o_1
XANTENNA__09063__B1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09366__B2 _04604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10144__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout304 _05458_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__buf_2
Xfanout315 _02288_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07377__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout326 net327 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_4
Xfanout337 _02110_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09933__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09813_ total_design.core.ctrl.instruction\[9\] total_design.core.ctrl.instruction\[10\]
+ net556 vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__nand3b_2
Xfanout359 _05017_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout386_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ _04121_ _04966_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__nor2_1
X_06956_ total_design.core.regFile.register\[11\]\[8\] net614 net595 total_design.core.regFile.register\[8\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__a22o_1
XANTENNA__12122__B1 _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13752__Q total_design.core.data_bus_o\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09675_ net313 net297 _04354_ _04900_ net289 vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__o32a_1
X_06887_ net752 _02442_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[6\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout553_A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06577__B net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08626_ total_design.lcd_display.cnt_500hz\[0\] net711 vssd1 vssd1 vccd1 vccd1 _00005_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_55_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06352__A1 total_design.core.ctrl.instruction\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_167_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ total_design.data_in_BUS\[13\] net342 _03903_ vssd1 vssd1 vccd1 vccd1 _03904_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_46_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08792__B _02515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07508_ total_design.core.regFile.register\[25\]\[18\] net842 net763 total_design.core.regFile.register\[6\]\[18\]
+ _03017_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__a221o_1
X_08488_ _03839_ _03840_ _03768_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07301__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07439_ total_design.core.regFile.register\[20\]\[17\] net670 net612 total_design.core.regFile.register\[11\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__a22o_1
XANTENNA__06655__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10319__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout606_X net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10450_ net199 net2437 net383 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07201__B _02718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09109_ net322 _04149_ net316 vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10381_ net212 net2608 net486 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12120_ total_design.lcd_display.row_2\[70\] _05819_ _05839_ total_design.lcd_display.row_1\[62\]
+ _05975_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12051_ _05801_ _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__nor2_1
XANTENNA__10054__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold380 total_design.lcd_display.row_2\[60\] vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold391 net98 vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11002_ _05257_ _05258_ _05260_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07907__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09843__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09109__A1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 _01945_ vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__buf_4
Xfanout871 net872 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_4
Xfanout882 net883 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__buf_2
Xfanout893 _02022_ vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__clkbuf_2
X_12953_ clknet_leaf_195_clk _00420_ net1009 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1080 total_design.core.regFile.register\[29\]\[7\] vssd1 vssd1 vccd1 vccd1 net2396
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08332__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1091 total_design.core.regFile.register\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 net2407
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ total_design.keypad0.key_out\[1\] total_design.keypad0.key_out\[3\] total_design.keypad0.key_out\[2\]
+ total_design.data_from_keypad\[0\] vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_107_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ clknet_leaf_141_clk _00351_ net1182 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07540__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11835_ total_design.lcd_display.currentState\[0\] total_design.lcd_display.currentState\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11613__S net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14554_ net1274 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XFILLER_0_135_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11766_ _01808_ _05693_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__nor2_2
XANTENNA__09293__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10737__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ clknet_leaf_122_clk _00972_ net1168 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14493__Q total_design.core.ctrl.instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10717_ net186 net2231 net359 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__mux2_1
XANTENNA__06646__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14485_ clknet_leaf_36_clk _01552_ net1072 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ net32 net936 _05690_ net1866 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13436_ clknet_leaf_30_clk _00903_ net1064 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10648_ net197 net2591 net477 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13367_ clknet_leaf_164_clk _00834_ net1164 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12444__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10579_ net211 net2112 net371 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12318_ net990 _01583_ _01584_ _01585_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07071__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13298_ clknet_leaf_145_clk _00765_ net1183 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12249_ _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07359__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09753__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06810_ total_design.core.regFile.register\[19\]\[5\] net825 net778 total_design.core.regFile.register\[22\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07790_ total_design.core.regFile.register\[11\]\[24\] net795 _03294_ _03295_ vssd1
+ vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__a211o_1
XANTENNA__12104__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08596__C net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06741_ total_design.core.regFile.register\[12\]\[4\] _01980_ net759 total_design.core.regFile.register\[21\]\[4\]
+ _02304_ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__a221o_1
X_09460_ total_design.core.math.pc_val\[18\] _04676_ vssd1 vssd1 vccd1 vccd1 _04696_
+ sky130_fd_sc_hd__xnor2_1
X_06672_ net333 net323 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__xnor2_4
XANTENNA__07531__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08411_ _01888_ _03719_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__nand2_2
X_09391_ net318 _04435_ _04629_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08342_ net1487 net939 _03705_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[28\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08273_ net1362 net560 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[23\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_129_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10139__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06637__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout134_A _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09928__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07224_ total_design.core.regFile.register\[20\]\[13\] net670 _02757_ _02759_ net686
+ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06563__D net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07155_ _02025_ _02695_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[11\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09587__B2 _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1043_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10197__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07086_ _02617_ _02626_ _02628_ _02630_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__or4_1
XANTENNA__07062__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09229__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13747__Q total_design.core.data_bus_o\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1210_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout134 _05686_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_2
Xfanout145 net146 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout670_A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout156 _05681_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08787__B total_design.core.data_mem.data_cpu_i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout167 net168 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout178 net179 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10602__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout189 net192 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_2
X_07988_ total_design.core.regFile.register\[0\]\[28\] net875 _03469_ _03485_ vssd1
+ vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__o22ai_4
XANTENNA__07036__X total_design.core.data_mem.data_cpu_i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ net168 net2078 net456 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06939_ _02449_ _02491_ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__xor2_4
XANTENNA_clkbuf_leaf_200_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08314__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09658_ _04874_ _04882_ _04884_ net450 vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ net1839 net338 net714 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[30\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__06876__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ total_design.core.math.pc_val\[24\] _04799_ vssd1 vssd1 vccd1 vccd1 _04819_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11620_ _05477_ net1718 net134 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__mux2_1
XANTENNA__09275__B1 _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11551_ net1770 _05651_ net146 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__mux2_1
XANTENNA__06628__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10049__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09838__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10502_ net261 net2310 net483 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__mux2_1
XANTENNA__06473__D net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14270_ clknet_leaf_47_clk _00002_ net1098 vssd1 vssd1 vccd1 vccd1 wishbone.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09027__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11482_ net1547 _05646_ net155 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__mux2_1
X_13221_ clknet_leaf_117_clk _00688_ net1161 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_150_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10433_ net257 net2309 net382 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07589__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ clknet_leaf_201_clk _00619_ net1004 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10364_ net276 net2561 net484 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12103_ total_design.lcd_display.row_1\[21\] _05826_ _05843_ total_design.lcd_display.row_1\[125\]
+ _05959_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_59_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ clknet_leaf_149_clk _00550_ net1148 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06800__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10295_ _04113_ _04968_ _05002_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__or3_1
X_12034_ net2883 _05847_ _05848_ total_design.lcd_display.row_2\[122\] _05893_ vssd1
+ vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__a221o_1
XANTENNA__11608__S net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09750__A1 total_design.core.regFile.register\[29\]\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10512__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13985_ clknet_leaf_96_clk _01165_ net1253 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08305__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12936_ clknet_leaf_169_clk _00403_ net1160 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09161__X _04409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_8__f_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ clknet_leaf_8_clk _00334_ net1016 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06867__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12439__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11818_ total_design.lcd_display.cnt_20ms\[10\] _05709_ net1858 vssd1 vssd1 vccd1
+ vccd1 _05712_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_174_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12798_ clknet_leaf_180_clk _00265_ net1044 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ net1309 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XANTENNA__11073__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11749_ net2866 net960 net293 total_design.core.data_bus_o\[21\] vssd1 vssd1 vccd1
+ vccd1 _01377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09748__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14468_ clknet_leaf_54_clk net1377 net1110 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07292__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13419_ clknet_leaf_120_clk _00886_ net1191 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07029__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07776__B _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14399_ clknet_leaf_44_clk _01536_ net1085 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08960_ _04212_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07911_ total_design.core.regFile.register\[7\]\[26\] net653 net605 total_design.core.regFile.register\[15\]\[26\]
+ _03411_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__a221o_1
X_08891_ _04143_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__and2b_1
XANTENNA__11518__S net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07842_ total_design.core.regFile.register\[25\]\[25\] net843 net832 total_design.core.regFile.register\[31\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__a22o_1
XANTENNA__10422__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07752__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07773_ _03254_ _03279_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__nand2_1
X_09512_ _04742_ _04744_ net707 vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__o21a_1
X_06724_ _02286_ net315 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__nand2_1
XANTENNA__06558__D net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11150__B1_N _05358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07504__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09443_ net903 _04678_ _04679_ _02346_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__o211ai_4
X_06655_ total_design.core.regFile.register\[30\]\[2\] net659 net569 total_design.core.regFile.register\[17\]\[2\]
+ _02222_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__a221o_1
XANTENNA__06858__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09257__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09374_ total_design.core.data_cpu_o\[14\] net756 _04608_ _04613_ vssd1 vssd1 vccd1
+ vccd1 _04614_ sky130_fd_sc_hd__a211o_1
X_06586_ total_design.core.regFile.register\[23\]\[1\] net746 net735 net732 vssd1
+ vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__and4_1
XFILLER_0_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08325_ total_design.core.data_mem.data_write_adr_reg\[20\] net546 net538 total_design.core.data_mem.data_read_adr_reg\[20\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout137_X net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08256_ net1317 net560 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[6\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_6_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07283__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07207_ _02689_ _02744_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__nor2_2
XFILLER_0_43_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08187_ net891 _03602_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[30\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11367__A1 _05411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1046_X net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_104_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07138_ total_design.core.regFile.register\[3\]\[11\] net866 net819 total_design.core.regFile.register\[17\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07440__C1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07069_ total_design.core.regFile.register\[18\]\[10\] net857 net798 total_design.core.regFile.register\[29\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07991__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ net183 net2114 net407 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10332__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_X net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13770_ clknet_leaf_55_clk total_design.core.data_mem.stored_data_adr\[13\] net1114
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_adr_o\[13\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12095__A2 _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ _05056_ _05170_ _05204_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__and3_1
X_12721_ clknet_leaf_150_clk _00188_ net1145 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_154_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06849__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11390__C _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12652_ clknet_leaf_118_clk _00119_ net1160 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06257__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09248__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06484__C net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11603_ _05671_ net1659 net138 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ clknet_leaf_176_clk _00050_ net1047 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14322_ clknet_leaf_68_clk _01483_ net1109 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_leaf_169_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire310 _02632_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_4
XFILLER_0_108_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11534_ net1571 _05679_ net147 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__mux2_1
XANTENNA__06781__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07274__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_122_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11399__A _05361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14253_ clknet_leaf_106_clk _01433_ net1234 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11465_ net1608 _05667_ net154 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__mux2_1
XANTENNA__10507__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13204_ clknet_leaf_141_clk _00671_ net1175 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10416_ net203 net1972 net387 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__mux2_1
XANTENNA__07026__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14184_ clknet_leaf_79_clk net1786 net1218 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11396_ net303 _05653_ _05654_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_78_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13135_ clknet_leaf_146_clk _00602_ net1178 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10347_ net218 net2244 net488 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07982__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13066_ clknet_leaf_19_clk _00533_ net1049 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10278_ net225 net2824 net499 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__mux2_1
XANTENNA__10750__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12017_ total_design.lcd_display.row_2\[105\] _05834_ _05841_ total_design.lcd_display.row_1\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10242__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06537__A1 total_design.core.ctrl.imm_32\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07734__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12086__A2 _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13968_ clknet_leaf_110_clk _01148_ net1225 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12919_ clknet_leaf_164_clk _00386_ net1164 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13899_ clknet_leaf_88_clk _01079_ net1260 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06440_ net971 _01916_ _02012_ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__nand3_1
XFILLER_0_174_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06394__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06371_ _01931_ net918 net928 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__and3b_4
XFILLER_0_145_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08890__B _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08110_ net750 _03602_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[30\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09090_ net463 _04242_ net328 vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08041_ total_design.core.regFile.register\[5\]\[29\] net628 net624 total_design.core.regFile.register\[14\]\[29\]
+ _03535_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10417__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold902 total_design.core.regFile.register\[15\]\[29\] vssd1 vssd1 vccd1 vccd1 net2218
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold913 total_design.core.regFile.register\[0\]\[13\] vssd1 vssd1 vccd1 vccd1 net2229
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12010__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold924 total_design.core.regFile.register\[31\]\[10\] vssd1 vssd1 vccd1 vccd1 net2240
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 total_design.core.regFile.register\[18\]\[2\] vssd1 vssd1 vccd1 vccd1 net2251
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 total_design.core.regFile.register\[14\]\[7\] vssd1 vssd1 vccd1 vccd1 net2262
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 total_design.core.regFile.register\[23\]\[25\] vssd1 vssd1 vccd1 vccd1 net2273
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08765__A2 _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold968 total_design.core.regFile.register\[16\]\[19\] vssd1 vssd1 vccd1 vccd1 net2284
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ net273 net2805 net417 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__mux2_1
Xhold979 total_design.core.regFile.register\[9\]\[9\] vssd1 vssd1 vccd1 vccd1 net2295
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06776__A1 _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07973__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08943_ net317 _04127_ _04193_ _04190_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__a31o_1
XANTENNA__08411__A _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10152__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08874_ net322 net312 _04104_ _04126_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_32_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11521__A1 _05477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1006_A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ _03329_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout466_A _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07756_ total_design.core.regFile.register\[13\]\[23\] net666 net636 total_design.core.regFile.register\[2\]\[23\]
+ _03262_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__a221o_1
XANTENNA__12077__A2 _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06707_ total_design.core.regFile.register\[9\]\[3\] net664 net567 total_design.core.regFile.register\[12\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a22o_1
XANTENNA__07489__C1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07687_ total_design.core.regFile.register\[25\]\[22\] net843 net765 total_design.core.regFile.register\[6\]\[22\]
+ _03196_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout633_A _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09426_ net701 _04661_ _04662_ _04105_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__o211a_1
X_06638_ total_design.core.regFile.register\[26\]\[2\] net869 net834 total_design.core.regFile.register\[10\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07968__Y _03467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09357_ _04549_ _04596_ net460 vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout800_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06569_ _02138_ _02139_ _02140_ _02141_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1163_X net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08308_ net1510 net940 _03688_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[11\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07697__A _03206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09288_ _04332_ _04529_ net319 vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08239_ net1378 net543 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[22\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__10327__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12537__B1 _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250_ _05414_ _05415_ _05417_ _05506_ _05507_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07008__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12001__A2 _05814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09402__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10201_ _04495_ net392 _04997_ vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_56_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11181_ net513 _05252_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__nand2_2
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10132_ net240 net1931 net399 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07208__Y _02746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ net251 net2573 net408 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__mux2_1
XANTENNA__10062__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11512__A1 _05648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09851__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11953__Y _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06479__C net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08975__B _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13822_ clknet_leaf_112_clk total_design.core.data_mem.data_cpu_i\[31\] net1207 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[31\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12068__A2 _05814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13753_ clknet_leaf_73_clk total_design.core.data_mem.stored_write_data\[28\] net1209
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[28\] sky130_fd_sc_hd__dfrtp_4
X_10965_ _05223_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08141__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12704_ clknet_leaf_1_clk _00171_ net1004 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13684_ clknet_leaf_50_clk total_design.core.data_mem.data_read_adr_i\[24\] net1097
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10896_ net520 _05154_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__nand2_2
XFILLER_0_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12635_ clknet_leaf_150_clk _00102_ net1147 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11621__S net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12566_ net1441 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07247__A2 _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10745__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11517_ net1849 _05650_ net151 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__mux2_1
X_14305_ clknet_leaf_104_clk _00019_ net1235 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10237__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12497_ net977 total_design.core.instr_mem.instruction_i\[12\] vssd1 vssd1 vccd1
+ vccd1 _01703_ sky130_fd_sc_hd__and2b_1
XFILLER_0_151_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12528__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14236_ clknet_leaf_57_clk _01416_ net1119 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dfrtp_1
Xhold209 net127 vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output95_A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11448_ net1695 _05645_ net157 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_169_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12452__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14167_ clknet_leaf_31_clk _01347_ net1061 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11379_ _05477_ _05624_ _05626_ _05637_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__and4_1
XANTENNA__11751__B2 total_design.core.data_bus_o\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13118_ clknet_leaf_157_clk _00585_ net1141 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14098_ clknet_leaf_86_clk _01278_ net1247 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_13049_ clknet_leaf_191_clk _00516_ net1012 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11503__A1 _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07707__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1260 net1261 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09761__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06389__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08885__B _02564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07610_ total_design.core.regFile.register\[19\]\[20\] net823 net810 total_design.core.regFile.register\[23\]\[20\]
+ _03115_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__a221o_1
XANTENNA__12059__A2 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08590_ _03895_ net880 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[11\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10700__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_clk sky130_fd_sc_hd__clkbuf_8
X_07541_ total_design.core.regFile.register\[20\]\[19\] net671 net634 total_design.core.regFile.register\[16\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__a22o_1
XANTENNA__13799__RESET_B net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07486__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07472_ total_design.core.ctrl.instruction\[18\] _02945_ vssd1 vssd1 vccd1 vccd1
+ _02994_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09211_ _02540_ net706 _04456_ _04105_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06423_ net928 net910 net907 vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09142_ _04215_ _04390_ net327 vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__mux2_1
XANTENNA__07238__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06354_ net966 net965 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__or2_1
XANTENNA__09632__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09073_ _04273_ _04249_ net467 vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__mux2_1
X_06285_ total_design.core.instr_mem.instruction_adr_i\[7\] total_design.core.instr_mem.instruction_adr_stored\[7\]
+ net984 vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10147__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout214_A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08024_ total_design.core.regFile.register\[29\]\[29\] net798 net763 total_design.core.regFile.register\[6\]\[29\]
+ _03519_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__a221o_1
XANTENNA__09936__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold710 total_design.core.regFile.register\[5\]\[2\] vssd1 vssd1 vccd1 vccd1 net2026
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold721 total_design.core.regFile.register\[16\]\[1\] vssd1 vssd1 vccd1 vccd1 net2037
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold732 total_design.core.regFile.register\[15\]\[13\] vssd1 vssd1 vccd1 vccd1 net2048
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11767__A net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold743 total_design.core.regFile.register\[31\]\[13\] vssd1 vssd1 vccd1 vccd1 net2059
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 total_design.core.regFile.register\[12\]\[20\] vssd1 vssd1 vccd1 vccd1 net2070
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1123_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold765 total_design.core.regFile.register\[12\]\[26\] vssd1 vssd1 vccd1 vccd1 net2081
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 total_design.core.regFile.register\[7\]\[22\] vssd1 vssd1 vccd1 vccd1 net2092
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11742__B2 total_design.core.data_bus_o\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold787 total_design.core.regFile.register\[31\]\[28\] vssd1 vssd1 vccd1 vccd1 net2103
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ net195 net2410 net418 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__mux2_1
Xhold798 total_design.core.regFile.register\[20\]\[26\] vssd1 vssd1 vccd1 vccd1 net2114
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07410__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13755__Q total_design.core.data_bus_o\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout583_A _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08926_ _03016_ _03064_ net470 vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09699__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1410 total_design.core.regFile.register\[11\]\[21\] vssd1 vssd1 vccd1 vccd1 net2726
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1421 total_design.core.regFile.register\[12\]\[9\] vssd1 vssd1 vccd1 vccd1 net2737
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1432 total_design.core.regFile.register\[17\]\[29\] vssd1 vssd1 vccd1 vccd1 net2748
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08857_ _01921_ _02014_ net888 net756 vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout750_A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1443 total_design.core.regFile.register\[12\]\[10\] vssd1 vssd1 vccd1 vccd1 net2759
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1454 total_design.core.regFile.register\[22\]\[22\] vssd1 vssd1 vccd1 vccd1 net2770
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout848_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1465 total_design.core.regFile.register\[15\]\[9\] vssd1 vssd1 vccd1 vccd1 net2781
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07808_ total_design.core.regFile.register\[2\]\[24\] net637 net605 total_design.core.regFile.register\[15\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__a22o_1
XANTENNA__08910__A2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1476 total_design.core.regFile.register\[21\]\[20\] vssd1 vssd1 vccd1 vccd1 net2792
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10610__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1487 total_design.core.regFile.register\[3\]\[3\] vssd1 vssd1 vccd1 vccd1 net2803
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08788_ _02666_ net300 vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_140_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1498 total_design.core.regFile.register\[12\]\[16\] vssd1 vssd1 vccd1 vccd1 net2814
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07739_ total_design.core.regFile.register\[24\]\[23\] net790 net758 total_design.core.regFile.register\[4\]\[23\]
+ _03246_ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10750_ net2875 net355 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_49_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07477__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09409_ _04461_ _04646_ net317 vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__mux2_1
XANTENNA__06685__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10681_ net197 net2299 net362 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout803_X net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11441__S net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12420_ _01674_ _01675_ _01676_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__a21o_1
XFILLER_0_168_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07229__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_7__f_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_97_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12351_ total_design.core.math.pc_val\[23\] net988 vssd1 vssd1 vccd1 vccd1 _01615_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10057__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11302_ _05521_ _05556_ _05558_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09846__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11948__Y _05810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12282_ total_design.core.math.pc_val\[15\] net524 _06120_ _06121_ vssd1 vssd1 vccd1
+ vccd1 _01485_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14021_ clknet_leaf_89_clk _01201_ net1258 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[103\]
+ sky130_fd_sc_hd__dfrtp_1
X_11233_ _05489_ _05491_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09418__Y _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11733__B2 total_design.core.data_bus_o\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11164_ net514 _05184_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__nand2_1
XANTENNA__06270__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07401__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ net173 total_design.core.regFile.register\[19\]\[28\] net404 vssd1 vssd1
+ vccd1 vccd1 _00419_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_164_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11095_ _01855_ _05024_ _05027_ _05353_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__and4_1
X_10046_ net184 net2852 net411 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_160_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold70 total_design.core.data_mem.data_cpu_i_reg\[9\] vssd1 vssd1 vccd1 vccd1 net1386
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11616__S net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 total_design.core.instr_mem.instruction_adr_stored\[4\] vssd1 vssd1 vccd1
+ vccd1 net1397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 total_design.core.math.pc_val\[20\] vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10520__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14496__Q total_design.core.ctrl.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13805_ clknet_leaf_76_clk total_design.core.data_mem.data_cpu_i\[14\] net1214 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[14\] sky130_fd_sc_hd__dfrtp_1
X_11997_ total_design.lcd_display.row_1\[72\] _05816_ _05841_ total_design.lcd_display.row_1\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a22o_1
XANTENNA__08114__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10948_ _05150_ _05175_ _05203_ _05205_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__a22o_1
X_13736_ clknet_leaf_76_clk total_design.core.data_mem.stored_write_data\[11\] net1214
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_133_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09862__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13667_ clknet_leaf_60_clk total_design.core.data_mem.data_read_adr_i\[7\] net1131
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[7\] sky130_fd_sc_hd__dfrtp_1
X_10879_ _05134_ _05136_ _05131_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__or3b_1
XANTENNA__12447__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12618_ clknet_leaf_21_clk _00085_ net1049 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13598_ clknet_leaf_61_clk net1320 net1129 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12549_ net1418 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06391__D net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09756__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 _01947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07640__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14219_ clknet_leaf_59_clk _01399_ net1126 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12774__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07928__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09393__A2 _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout508 _04103_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__buf_4
Xfanout519 _01886_ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06600__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09760_ net237 net2352 net442 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__mux2_1
X_06972_ total_design.core.regFile.register\[9\]\[8\] net852 net821 total_design.core.regFile.register\[17\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__a22o_1
X_08711_ total_design.keypad0.counter\[6\] _03952_ total_design.keypad0.counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__a21oi_1
X_09691_ _03553_ _04186_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__nand2_1
XANTENNA__11526__S net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1090 net1096 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09063__Y _04315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08642_ net712 _03928_ _03929_ _03930_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__and4_1
XANTENNA__10430__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06364__C1 total_design.core.ctrl.instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_174_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08573_ net1739 net342 net720 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[28\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_77_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07524_ _03041_ _03042_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__nand2_1
XANTENNA__07459__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11660__A0 _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07455_ total_design.core.regFile.register\[3\]\[17\] net865 net819 total_design.core.regFile.register\[17\]\[17\]
+ _02970_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout331_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06406_ net925 net919 net914 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__and3_1
XFILLER_0_174_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09605__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07386_ total_design.core.regFile.register\[31\]\[16\] net603 net595 total_design.core.regFile.register\[8\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06582__C net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09125_ net281 net2044 net453 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__mux2_1
XANTENNA__10215__A1 _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06337_ wishbone.curr_state\[2\] _01731_ _01907_ wishbone.curr_state\[0\] vssd1 vssd1
+ vccd1 vccd1 _00002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1240_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09056_ net459 _04152_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__nand2_1
X_06268_ total_design.core.data_adr_o\[24\] _01846_ net961 vssd1 vssd1 vccd1 vccd1
+ _01847_ sky130_fd_sc_hd__mux2_2
XANTENNA__07631__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout798_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ total_design.core.regFile.register\[10\]\[28\] net617 _03503_ net687 vssd1
+ vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_92_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold540 total_design.lcd_display.row_2\[98\] vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10605__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06199_ net1799 _01761_ _01778_ vssd1 vssd1 vccd1 vccd1 total_design.core.mem_ctrl.next_state\[1\]
+ sky130_fd_sc_hd__a21oi_1
Xhold551 total_design.core.math.pc_val\[24\] vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 total_design.lcd_display.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 total_design.core.regFile.register\[30\]\[1\] vssd1 vssd1 vccd1 vccd1 net1889
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 total_design.core.regFile.register\[31\]\[2\] vssd1 vssd1 vccd1 vccd1 net1900
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold595 total_design.core.regFile.register\[15\]\[4\] vssd1 vssd1 vccd1 vccd1 net1911
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout586_X net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15__f_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_70_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09958_ net272 net2058 net420 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ net471 _03595_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__A1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13862__D total_design.core.ctrl.imm_32\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ net260 net2624 net427 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__mux2_1
Xhold1240 total_design.core.regFile.register\[18\]\[12\] vssd1 vssd1 vccd1 vccd1 net2556
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 total_design.core.regFile.register\[18\]\[16\] vssd1 vssd1 vccd1 vccd1 net2567
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ _05795_ total_design.keypad0.key_out\[2\] net530 vssd1 vssd1 vccd1 vccd1
+ _01449_ sky130_fd_sc_hd__mux2_1
Xhold1262 total_design.core.regFile.register\[13\]\[30\] vssd1 vssd1 vccd1 vccd1 net2578
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10340__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07698__A2 _03206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1273 total_design.core.regFile.register\[20\]\[14\] vssd1 vssd1 vccd1 vccd1 net2589
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1284 total_design.core.regFile.register\[15\]\[31\] vssd1 vssd1 vccd1 vccd1 net2600
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1295 total_design.core.regFile.register\[5\]\[20\] vssd1 vssd1 vccd1 vccd1 net2611
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11851_ total_design.lcd_display.currentState\[0\] _05719_ _05728_ _05736_ vssd1
+ vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_68_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ net517 _05059_ _05060_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_68_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11782_ net1656 net954 _05699_ _01784_ vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11651__A0 _05630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13521_ clknet_leaf_152_clk _00988_ net1146 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10733_ total_design.core.regFile.register\[0\]\[8\] net356 vssd1 vssd1 vccd1 vccd1
+ _01007_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ clknet_leaf_169_clk _00919_ net1160 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10664_ net258 net2075 net363 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12403_ net992 _04907_ net894 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13383_ clknet_leaf_176_clk _00850_ net1052 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10595_ net277 net2222 net366 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12334_ _01596_ _01598_ _01595_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07083__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06830__B1 _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12265_ net902 _02845_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10515__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14004_ clknet_leaf_99_clk _01184_ net1227 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11216_ _05473_ _05474_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__nand2_1
XANTENNA__08032__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12196_ _06043_ _06044_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__nor2_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__clkbuf_4
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__clkbuf_4
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__clkbuf_4
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__clkbuf_4
X_11147_ _05358_ _05405_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11078_ net351 _05155_ _05328_ _05330_ _05336_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__o2111a_1
XANTENNA__10250__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ net249 net2483 net412 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__mux2_1
XANTENNA__07689__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06897__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06386__D net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11642__A0 _05612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06649__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13719_ clknet_leaf_34_clk total_design.core.data_mem.stored_read_data\[26\] net1067
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07240_ total_design.core.regFile.register\[31\]\[13\] net831 net806 total_design.core.regFile.register\[5\]\[13\]
+ _02775_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07861__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07171_ total_design.core.regFile.register\[13\]\[12\] net669 net565 total_design.core.regFile.register\[3\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07074__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07613__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06821__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10425__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09366__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout316 net317 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_2
X_09812_ net163 net2752 net439 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__mux2_1
Xfanout327 _02236_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_4
Xfanout338 net343 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06955_ total_design.core.regFile.register\[15\]\[8\] net606 net584 total_design.core.regFile.register\[6\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__a22o_1
X_09743_ net905 _04964_ _04965_ _04963_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__o211a_4
XANTENNA_fanout281_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10160__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09674_ _04812_ _04899_ net330 vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__mux2_1
X_06886_ _02399_ _02441_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__xor2_2
X_08625_ _03912_ _03914_ _03915_ _03916_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__nor4_1
XANTENNA_fanout1190_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06352__A2 total_design.core.ctrl.instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A total_design.core.data_mem.next_write vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_89_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08556_ _03899_ _03902_ _03768_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_46_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11633__A0 _05679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07507_ _03022_ _03024_ _03026_ _03027_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__or4_1
XFILLER_0_92_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08487_ _03817_ _03819_ _03838_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07438_ _02956_ _02958_ _02960_ _02961_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07852__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07369_ total_design.core.ctrl.instruction\[28\] net889 vssd1 vssd1 vccd1 vccd1 _02897_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout501_X net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09108_ net324 _04141_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__nor2_1
XANTENNA__07065__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380_ net218 net2621 net484 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__mux2_1
XANTENNA__07604__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09039_ _02238_ net448 net289 _04290_ _04286_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__o221a_1
XFILLER_0_62_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10335__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12050_ _05754_ _05817_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold370 total_design.lcd_display.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 total_design.lcd_display.row_2\[29\] vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_X net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold392 _01359_ vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ _05231_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout968_X net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout850 _01951_ vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_8
Xfanout861 net864 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09425__A _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout872 _01938_ vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__buf_4
XFILLER_0_99_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout883 _03671_ vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__clkbuf_4
Xfanout894 net895 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__buf_2
XANTENNA__10070__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12952_ clknet_leaf_138_clk _00419_ net1184 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1070 total_design.core.regFile.register\[20\]\[28\] vssd1 vssd1 vccd1 vccd1 net2386
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 total_design.core.regFile.register\[8\]\[24\] vssd1 vssd1 vccd1 vccd1 net2397
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06487__C net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11903_ total_design.keypad0.key_counter\[1\] total_design.keypad0.key_counter\[0\]
+ total_design.keypad0.key_counter\[2\] total_design.keypad0.key_counter\[3\] vssd1
+ vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__and4_1
XANTENNA__11961__Y _05823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1092 total_design.core.regFile.register\[10\]\[31\] vssd1 vssd1 vccd1 vccd1 net2408
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ clknet_leaf_178_clk _00350_ net1033 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _05719_ _05720_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__nand2_1
XANTENNA__06784__A total_design.core.ctrl.instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09160__A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14553_ net1273 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
X_11765_ net1809 net956 _05698_ _01858_ vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08096__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ clknet_leaf_201_clk _00971_ net1003 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10716_ net189 net2307 net360 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__mux2_1
X_11696_ net31 net935 net878 net1825 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__o22a_1
X_14484_ clknet_leaf_37_clk _01551_ net1077 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07843__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13435_ clknet_leaf_147_clk _00902_ net1152 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10647_ net202 net2398 net477 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07056__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13366_ clknet_leaf_154_clk _00833_ net1136 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10578_ net217 net2677 net369 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__mux2_1
XANTENNA__10753__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14201__RESET_B net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06803__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12317_ net990 _04717_ net894 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10245__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13297_ clknet_leaf_151_clk _00764_ net1145 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12248_ total_design.core.math.pc_val\[12\] total_design.core.program_count.imm_val_reg\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12179_ _06020_ _06022_ _06027_ _06028_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__o211a_1
XANTENNA__08020__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12460__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06740_ total_design.core.regFile.register\[9\]\[4\] net850 net819 total_design.core.regFile.register\[17\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06397__C _01950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06671_ net333 net332 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__nand2_1
XANTENNA__08893__B _02367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ _03745_ _03765_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09390_ net314 _04433_ net296 vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11615__A0 _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08341_ total_design.core.data_mem.data_write_adr_reg\[28\] net547 net539 total_design.core.data_mem.data_read_adr_reg\[28\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08087__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11105__A total_design.core.data_bus_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08272_ net1374 net557 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[22\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07295__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07834__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07223_ total_design.core.regFile.register\[21\]\[13\] net597 net589 total_design.core.regFile.register\[1\]\[13\]
+ _02758_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12477__A_N net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07154_ total_design.core.ctrl.instruction\[5\] _02694_ vssd1 vssd1 vccd1 vccd1 _02695_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA__12040__B1 _05850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07085_ total_design.core.regFile.register\[30\]\[10\] net838 net834 total_design.core.regFile.register\[10\]\[10\]
+ _02629_ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__a221o_1
XANTENNA__10155__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09229__B _04474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1036_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09944__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09339__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout496_A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout135 _05686_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1203_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout146 _05683_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 net158 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout168 _04950_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_1
X_07987_ _03474_ _03476_ _03478_ _03484_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__or4_1
Xfanout179 _04890_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout663_A _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06573__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06938_ _02489_ _02490_ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__nand2_2
X_09726_ net507 _04949_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_87_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09657_ _03462_ net448 _04879_ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__o211a_1
X_06869_ total_design.core.regFile.register\[9\]\[6\] net852 net829 total_design.core.regFile.register\[1\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout451_X net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08608_ total_design.data_in_BUS\[29\] net341 net715 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[29\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_139_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09588_ _04810_ _04814_ _04817_ net450 vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__a31o_1
XANTENNA__11606__A0 _05652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08539_ _03876_ _03885_ _03887_ _03886_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__a31o_1
XANTENNA__08078__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09275__B2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11550_ net1640 _05650_ net148 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07286__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10501_ net267 net2247 net481 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11481_ net1684 _05645_ net153 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__mux2_1
XANTENNA__09027__A1 total_design.core.math.pc_val\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ clknet_leaf_128_clk _00687_ net1194 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10432_ net280 net2452 net381 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__mux2_1
XANTENNA__12031__B1 _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13151_ clknet_leaf_181_clk _00618_ net1043 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10065__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10363_ net244 net2237 net485 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__mux2_1
XANTENNA__10593__A0 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12102_ total_design.lcd_display.row_2\[109\] _05834_ _05841_ total_design.lcd_display.row_1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09854__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11956__Y _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13082_ clknet_leaf_125_clk _00549_ net1189 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10294_ net161 net2416 net498 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__mux2_1
X_12033_ total_design.lcd_display.row_2\[106\] _05834_ _05852_ total_design.lcd_display.row_2\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__a22o_1
XANTENNA__08002__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06498__B net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 net681 vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__buf_4
Xfanout691 net694 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_8
X_13984_ clknet_leaf_110_clk _01164_ net1227 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12935_ clknet_leaf_175_clk _00402_ net1053 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11624__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12866_ clknet_leaf_131_clk _00333_ net1197 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10748__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08069__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11817_ total_design.lcd_display.cnt_20ms\[11\] total_design.lcd_display.cnt_20ms\[10\]
+ _05709_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_174_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ clknet_leaf_10_clk _00264_ net1019 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08218__B net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11073__A1 total_design.core.data_bus_o\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07277__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ net1308 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_172_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11748_ net1732 net958 net291 total_design.core.data_bus_o\[20\] vssd1 vssd1 vccd1
+ vccd1 _01376_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07816__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14467_ clknet_leaf_54_clk net1447 net1110 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12455__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11679_ _05645_ net1800 net129 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07029__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12022__B1 _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13418_ clknet_leaf_25_clk _00885_ net1106 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14398_ clknet_leaf_44_clk _01535_ net1085 vssd1 vssd1 vccd1 vccd1 total_design.keypad0.key_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13349_ clknet_leaf_116_clk _00816_ net1203 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09764__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07910_ total_design.core.regFile.register\[14\]\[26\] net625 net583 total_design.core.regFile.register\[6\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__a22o_1
XANTENNA__10703__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08890_ net334 _02468_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__or2_1
XANTENNA__09065__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07841_ total_design.core.regFile.register\[29\]\[25\] net799 net777 total_design.core.regFile.register\[22\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__a22o_1
XANTENNA__12089__B1 _05850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07772_ _03276_ _03277_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09511_ _03137_ _03185_ _04722_ _04743_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a31o_1
X_06723_ net551 _02263_ _02266_ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11534__S net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ total_design.core.data_cpu_o\[17\] net755 _04124_ _04675_ vssd1 vssd1 vccd1
+ vccd1 _04679_ sky130_fd_sc_hd__a22oi_2
X_06654_ total_design.core.regFile.register\[29\]\[2\] net658 net593 total_design.core.regFile.register\[8\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09373_ net967 net888 _04612_ net906 vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06585_ total_design.core.regFile.register\[15\]\[1\] net741 net732 net726 vssd1
+ vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_25_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08324_ net1490 net938 _03696_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[19\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09939__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07268__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12261__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07807__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08255_ net1473 net560 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[5\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout411_A net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07206_ _02587_ _02637_ _02638_ _02690_ _02634_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__o311a_1
XANTENNA__12013__B1 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08186_ net891 _03559_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[29\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06216__X _01795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06590__C net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07137_ total_design.core.regFile.register\[12\]\[11\] net774 net772 total_design.core.regFile.register\[28\]\[11\]
+ _02678_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07068_ _02598_ _02600_ _02612_ net682 total_design.core.regFile.register\[0\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__o32a_4
XTAP_TAPCELL_ROW_37_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout780_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06794__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11110__C_N _05028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10613__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout666_X net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06886__X _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09709_ _03598_ _03599_ _04932_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__a21oi_1
X_10981_ _05056_ _05239_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__nand2_1
XANTENNA__13870__D total_design.core.ctrl.imm_32\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout833_X net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11444__S net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12720_ clknet_leaf_184_clk _00187_ net1039 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12651_ clknet_leaf_127_clk _00118_ net1191 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11390__D _05648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_0__f_clk_X clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ _05680_ net1808 net140 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__mux2_1
XANTENNA__12252__B1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12582_ clknet_leaf_195_clk _00049_ net1008 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10802__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14321_ clknet_leaf_67_clk _01482_ net1111 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[12\]
+ sky130_fd_sc_hd__dfrtp_4
Xwire300 _02686_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11533_ net1526 _05632_ net146 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__mux2_1
Xwire311 _02418_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11464_ net1665 _05665_ net153 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__mux2_1
XANTENNA__12004__B1 _05834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14252_ clknet_leaf_106_clk _01432_ net1234 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13203_ clknet_leaf_190_clk _00670_ net1034 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10415_ net208 net2027 net385 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14183_ clknet_leaf_79_clk net1683 net1218 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
X_11395_ net513 _05054_ _05459_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_78_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13134_ clknet_leaf_188_clk _00601_ net1028 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10346_ net213 net2653 net488 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__mux2_1
XANTENNA__07431__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13065_ clknet_leaf_177_clk _00532_ net1047 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10523__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10277_ net233 net2016 net497 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12016_ total_design.lcd_display.row_1\[65\] _05804_ _05818_ total_design.lcd_display.row_2\[81\]
+ _05872_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__a221o_1
XANTENNA__14499__Q total_design.core.ctrl.instruction\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_174_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08931__B1 _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13967_ clknet_leaf_84_clk _01147_ net1247 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10759__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12918_ clknet_leaf_156_clk _00385_ net1142 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07498__B1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13898_ clknet_leaf_87_clk _01078_ net1250 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12849_ clknet_leaf_150_clk _00316_ net1147 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09759__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06370_ total_design.core.regFile.register\[18\]\[0\] net927 net949 net917 vssd1
+ vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__nand4_1
XFILLER_0_174_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14519_ net1291 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_56_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08040_ total_design.core.regFile.register\[20\]\[29\] net670 net569 total_design.core.regFile.register\[17\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold903 total_design.core.regFile.register\[7\]\[24\] vssd1 vssd1 vccd1 vccd1 net2219
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold914 total_design.core.regFile.register\[11\]\[22\] vssd1 vssd1 vccd1 vccd1 net2230
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 total_design.core.regFile.register\[19\]\[11\] vssd1 vssd1 vccd1 vccd1 net2241
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold936 total_design.core.regFile.register\[1\]\[8\] vssd1 vssd1 vccd1 vccd1 net2252
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08899__A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold947 total_design.keypad0.key_counter\[3\] vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09347__X _04588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold958 total_design.core.regFile.register\[22\]\[15\] vssd1 vssd1 vccd1 vccd1 net2274
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 total_design.core.regFile.register\[1\]\[10\] vssd1 vssd1 vccd1 vccd1 net2285
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ net257 net1978 net416 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__mux2_1
XANTENNA__11529__S net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06776__A2 total_design.core.data_mem.data_cpu_i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_11__f_clk_X clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ net320 _04193_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__nand2_1
XANTENNA__10433__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09175__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ net322 _04126_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__nor2_1
XANTENNA__06528__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14202__Q net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07824_ _03327_ _03328_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07755_ total_design.core.regFile.register\[26\]\[23\] net644 net562 total_design.core.regFile.register\[3\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout361_A net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06706_ total_design.core.regFile.register\[11\]\[3\] net613 net574 total_design.core.regFile.register\[24\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07686_ total_design.core.regFile.register\[31\]\[22\] net832 net777 total_design.core.regFile.register\[22\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07043__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06637_ total_design.core.regFile.register\[14\]\[2\] net864 net802 total_design.core.regFile.register\[8\]\[2\]
+ _02190_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__a221o_1
X_09425_ _02993_ net702 vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout247_X net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout626_A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12234__B1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06568_ total_design.core.regFile.register\[4\]\[1\] _02004_ _02122_ _02124_ _02137_
+ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__a2111o_1
X_09356_ _04129_ _04133_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08307_ total_design.core.data_mem.data_write_adr_reg\[11\] net548 net540 total_design.core.data_mem.data_read_adr_reg\[11\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__a221o_1
X_09287_ _04529_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10608__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06499_ total_design.core.regFile.register\[18\]\[0\] net747 net736 net730 vssd1
+ vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__and4_1
XFILLER_0_133_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08238_ net1442 net543 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[21\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07661__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout995_A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08169_ net892 _02746_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[12\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10200_ net2383 net392 vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_56_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11180_ _05357_ _05437_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_56_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13865__D total_design.core.ctrl.imm_32\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11439__S net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10131_ net254 net2648 net398 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10343__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10062_ net262 total_design.core.regFile.register\[20\]\[8\] net408 vssd1 vssd1 vccd1
+ vccd1 _00367_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_145_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07177__C1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06479__D net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07192__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13821_ clknet_leaf_113_clk total_design.core.data_mem.data_cpu_i\[30\] net1206 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[30\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09469__A1 _03090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06268__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13752_ clknet_leaf_72_clk total_design.core.data_mem.stored_write_data\[27\] net1205
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_74_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10964_ _05221_ _05222_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06495__C net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12703_ clknet_leaf_156_clk _00170_ net1140 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13683_ clknet_leaf_50_clk total_design.core.data_mem.data_read_adr_i\[23\] net1100
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[23\] sky130_fd_sc_hd__dfrtp_1
X_10895_ total_design.core.data_bus_o\[5\] net699 vssd1 vssd1 vccd1 vccd1 _05154_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12634_ clknet_leaf_134_clk _00101_ net1195 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12565_ net1448 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10518__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14304_ clknet_leaf_104_clk _00018_ net1235 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11516_ net1543 _05633_ net150 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__mux2_1
XANTENNA__07652__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12496_ net975 total_design.core.ctrl.instruction\[11\] net883 _01702_ vssd1 vssd1
+ vccd1 vccd1 _01550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14235_ clknet_leaf_57_clk _01415_ net1118 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11447_ net1561 _05643_ net157 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06207__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07404__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11378_ _05634_ _05635_ _05636_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14166_ clknet_leaf_32_clk _01346_ net1061 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06758__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13117_ clknet_leaf_11_clk _00584_ net1025 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10329_ net287 net1860 net491 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__mux2_1
XANTENNA__10253__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14097_ clknet_leaf_97_clk _01277_ net1246 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08231__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13048_ clknet_leaf_124_clk _00515_ net1186 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1250 net1251 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__clkbuf_4
Xfanout1261 net1264 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_1_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07183__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06930__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ total_design.core.regFile.register\[27\]\[19\] net578 net574 total_design.core.regFile.register\[24\]\[19\]
+ _03057_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__a221o_1
XFILLER_0_163_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07471_ net750 _02993_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[17\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09210_ net706 _04455_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__nand2_1
X_06422_ total_design.core.regFile.register\[6\]\[0\] net922 net917 net907 vssd1 vssd1
+ vccd1 vccd1 _01998_ sky130_fd_sc_hd__and4_1
XFILLER_0_158_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09141_ _04330_ _04389_ net461 vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06353_ net966 net965 vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__nor2_1
XANTENNA__10428__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09072_ _04321_ _04322_ net329 vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06284_ total_design.core.data_adr_o\[6\] _01862_ net964 vssd1 vssd1 vccd1 vccd1
+ _01863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08023_ total_design.core.regFile.register\[25\]\[29\] net842 net838 total_design.core.regFile.register\[30\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__a22o_1
XANTENNA__06997__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold700 total_design.core.regFile.register\[14\]\[14\] vssd1 vssd1 vccd1 vccd1 net2016
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout207_A _04740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold711 total_design.core.regFile.register\[10\]\[20\] vssd1 vssd1 vccd1 vccd1 net2027
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold722 total_design.core.regFile.register\[28\]\[5\] vssd1 vssd1 vccd1 vccd1 net2038
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 total_design.core.regFile.register\[14\]\[4\] vssd1 vssd1 vccd1 vccd1 net2049
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11767__B _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold744 total_design.core.regFile.register\[4\]\[11\] vssd1 vssd1 vccd1 vccd1 net2060
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold755 total_design.core.regFile.register\[17\]\[14\] vssd1 vssd1 vccd1 vccd1 net2071
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_153_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold766 total_design.core.regFile.register\[18\]\[18\] vssd1 vssd1 vccd1 vccd1 net2082
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 total_design.core.regFile.register\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 net2093
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 total_design.core.regFile.register\[16\]\[31\] vssd1 vssd1 vccd1 vccd1 net2104
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10163__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09974_ net198 net2122 net419 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__mux2_1
Xhold799 total_design.core.regFile.register\[3\]\[27\] vssd1 vssd1 vccd1 vccd1 net2115
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1116_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07038__A _02564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ _04175_ _04178_ net464 vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1400 total_design.core.regFile.register\[20\]\[5\] vssd1 vssd1 vccd1 vccd1 net2716
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout576_A _02089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1411 total_design.core.regFile.register\[22\]\[7\] vssd1 vssd1 vccd1 vccd1 net2727
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 total_design.core.regFile.register\[25\]\[11\] vssd1 vssd1 vccd1 vccd1 net2738
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 total_design.core.regFile.register\[29\]\[20\] vssd1 vssd1 vccd1 vccd1 net2749
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08856_ net972 _01918_ _04110_ net906 vssd1 vssd1 vccd1 vccd1 total_design.core.branch_ff
+ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_168_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07174__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1444 total_design.core.regFile.register\[30\]\[8\] vssd1 vssd1 vccd1 vccd1 net2760
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09253__A _02565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1455 total_design.core.regFile.register\[9\]\[29\] vssd1 vssd1 vccd1 vccd1 net2771
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07807_ total_design.core.regFile.register\[20\]\[24\] net671 net563 total_design.core.regFile.register\[3\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__a22o_1
Xhold1466 total_design.core.regFile.register\[5\]\[10\] vssd1 vssd1 vccd1 vccd1 net2782
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1477 total_design.core.regFile.register\[0\]\[14\] vssd1 vssd1 vccd1 vccd1 net2793
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08787_ _02770_ total_design.core.data_mem.data_cpu_i\[13\] vssd1 vssd1 vccd1 vccd1
+ _04042_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout743_A _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout364_X net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1488 total_design.core.regFile.register\[28\]\[8\] vssd1 vssd1 vccd1 vccd1 net2804
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06921__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 net128 vssd1 vssd1 vccd1 vccd1 net2815 sky130_fd_sc_hd__dlygate4sd3_1
X_07738_ total_design.core.regFile.register\[15\]\[23\] net846 _01980_ total_design.core.regFile.register\[12\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout910_A _01950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07669_ net553 _03157_ _03179_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_49_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09408_ _04550_ _04645_ net326 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__mux2_1
X_10680_ net201 net2717 net362 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__mux2_1
XANTENNA__07882__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09339_ _02795_ net508 net298 _04578_ _04579_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__o221a_1
XANTENNA__10338__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12350_ total_design.core.math.pc_val\[23\] net988 vssd1 vssd1 vccd1 vccd1 _01614_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11430__A1 _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07634__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout998_X net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11301_ _05556_ _05558_ _05521_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__a21oi_1
X_12281_ net900 _02893_ net524 vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11232_ _05389_ _05485_ _05486_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__and3_1
X_14020_ clknet_leaf_100_clk _01200_ net1228 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06404__X _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ _05420_ _05421_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__and2_1
XANTENNA__10073__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10114_ net178 net2133 net404 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__mux2_1
XANTENNA__09862__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11964__Y _05826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11094_ _05311_ _05320_ _05325_ _05352_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_164_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10045_ net187 net1949 net412 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__mux2_1
XANTENNA__06787__A _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07165__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 total_design.core.data_mem.data_cpu_i_reg\[21\] vssd1 vssd1 vccd1 vccd1 net1376
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 total_design.core.instr_mem.instruction_adr_stored\[5\] vssd1 vssd1 vccd1
+ vccd1 net1387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 total_design.core.instr_mem.instruction_adr_stored\[6\] vssd1 vssd1 vccd1
+ vccd1 net1398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 total_design.core.instr_mem.instruction_adr_stored\[19\] vssd1 vssd1 vccd1
+ vccd1 net1409 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output126_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06912__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13804_ clknet_leaf_76_clk total_design.core.data_mem.data_cpu_i\[13\] net1213 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11996_ total_design.lcd_display.row_1\[88\] _05812_ _05829_ total_design.lcd_display.row_1\[104\]
+ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__a22o_1
X_13735_ clknet_leaf_77_clk total_design.core.data_mem.stored_write_data\[10\] net1213
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[10\] sky130_fd_sc_hd__dfrtp_1
X_10947_ _05203_ _05205_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__nand2_1
XANTENNA__11632__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13666_ clknet_leaf_60_clk total_design.core.data_mem.data_read_adr_i\[6\] net1131
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[6\] sky130_fd_sc_hd__dfrtp_1
X_10878_ _05130_ _05136_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__nor2_1
XANTENNA__09102__S net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10756__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12617_ clknet_leaf_17_clk _00084_ net1046 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10248__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13597_ clknet_leaf_62_clk net1322 net1129 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08226__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11421__A1 _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12548_ net1468 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06979__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10772__A total_design.core.data_bus_o\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ net980 net2845 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__and2b_1
XANTENNA_2 _01999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__X _05479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14218_ clknet_leaf_59_clk _01398_ net1127 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14149_ clknet_leaf_43_clk _01329_ net1083 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08050__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout509 _04103_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_2
XANTENNA__09393__A3 _04631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09772__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06971_ total_design.core.regFile.register\[11\]\[8\] net796 net761 total_design.core.regFile.register\[21\]\[8\]
+ _02521_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08710_ _03971_ _00035_ _03974_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__nor3_2
XANTENNA__11488__A1 _05477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10711__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ _04912_ _04914_ _03559_ net707 vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06697__A _02263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1080 net1081 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__buf_2
Xfanout1091 net1096 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__clkbuf_2
X_08641_ total_design.lcd_display.cnt_500hz\[3\] _03921_ vssd1 vssd1 vccd1 vccd1 _03930_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06364__B1 total_design.core.ctrl.instruction\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__06903__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08572_ net1635 net342 net720 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[27\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__06984__X total_design.core.data_mem.data_cpu_i\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_53_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07523_ total_design.core.ctrl.instruction\[19\] _02994_ vssd1 vssd1 vccd1 vccd1
+ _03042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11542__S net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout157_A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07454_ total_design.core.regFile.register\[26\]\[17\] net869 net763 total_design.core.regFile.register\[6\]\[17\]
+ _02974_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07864__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06405_ _01739_ total_design.core.regFile.register\[12\]\[0\] net918 _01948_ vssd1
+ vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_79_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10158__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07385_ _02905_ _02907_ _02909_ _02911_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__or4_1
XFILLER_0_91_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06336_ wishbone.curr_state\[1\] _01731_ _01909_ wishbone.curr_state\[0\] vssd1 vssd1
+ vccd1 vccd1 _00001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09124_ _04370_ _04373_ net452 vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09947__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10215__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06582__D net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09055_ _04140_ _04145_ net459 vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__mux2_1
X_06267_ total_design.core.instr_mem.instruction_adr_i\[24\] total_design.core.instr_mem.instruction_adr_stored\[24\]
+ net982 vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08006_ total_design.core.regFile.register\[23\]\[28\] net679 net630 total_design.core.regFile.register\[5\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__a22o_1
Xhold530 total_design.lcd_display.row_2\[57\] vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06198_ total_design.core.mem_ctrl.state\[2\] _01764_ _01777_ vssd1 vssd1 vccd1 vccd1
+ _01778_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout693_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold541 total_design.data_in_BUS\[14\] vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold552 total_design.core.data_mem.data_bus_i_reg\[15\] vssd1 vssd1 vccd1 vccd1 net1868
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold563 total_design.lcd_display.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08041__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold574 total_design.core.regFile.register\[10\]\[16\] vssd1 vssd1 vccd1 vccd1 net1890
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold585 total_design.core.regFile.register\[29\]\[1\] vssd1 vssd1 vccd1 vccd1 net1901
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 total_design.core.regFile.register\[14\]\[27\] vssd1 vssd1 vccd1 vccd1 net1912
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07395__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09957_ net257 net2501 net420 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_X net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11479__A1 _05648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ _04160_ _04161_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__and2_1
XANTENNA__10621__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09888_ net281 net2455 net426 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__mux2_1
XANTENNA__07147__A2 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1230 total_design.core.regFile.register\[22\]\[4\] vssd1 vssd1 vccd1 vccd1 net2546
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12140__A2 _05830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09541__B1 _04410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1241 total_design.core.regFile.register\[24\]\[19\] vssd1 vssd1 vccd1 vccd1 net2557
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 total_design.core.regFile.register\[25\]\[9\] vssd1 vssd1 vccd1 vccd1 net2568
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ _04012_ _04093_ _04022_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__or3b_1
Xhold1263 total_design.core.regFile.register\[19\]\[15\] vssd1 vssd1 vccd1 vccd1 net2579
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09670__A2_N net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1274 total_design.core.regFile.register\[6\]\[18\] vssd1 vssd1 vccd1 vccd1 net2590
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1285 total_design.core.regFile.register\[20\]\[31\] vssd1 vssd1 vccd1 vccd1 net2601
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1296 total_design.keypad0.counter\[17\] vssd1 vssd1 vccd1 vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
X_11850_ _01724_ _05720_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__and2_1
X_10801_ total_design.core.data_bus_o\[11\] _01852_ _01884_ _05049_ vssd1 vssd1 vccd1
+ vccd1 _05060_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_68_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _01890_ _05693_ net953 net1778 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_67_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11452__S net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13520_ clknet_leaf_185_clk _00987_ net1037 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07855__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10732_ net2660 net354 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13451_ clknet_leaf_114_clk _00918_ net1204 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10663_ net281 net2365 net361 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__mux2_1
XANTENNA__10068__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12402_ _01658_ _01659_ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__or2_1
XANTENNA__09857__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11959__Y _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07607__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13382_ clknet_leaf_199_clk _00849_ net1001 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10594_ net246 net2348 net365 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11688__A total_design.bus_full vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12333_ _01595_ _01596_ _01598_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06281__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06830__A1 _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12264_ net2885 net525 _06104_ _06105_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14003_ clknet_leaf_92_clk _01183_ net1263 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11215_ _05461_ _05466_ _05451_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__o21ai_2
XANTENNA__08032__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12195_ total_design.core.math.pc_val\[6\] total_design.core.program_count.imm_val_reg\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__nor2_1
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__clkbuf_4
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07386__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__clkbuf_4
X_11146_ _05392_ _05400_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__xnor2_1
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
X_11077_ _05331_ _05334_ _05335_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__and3_1
XANTENNA__10531__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12131__A2 _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09532__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ net264 net2679 net412 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__mux2_1
XANTENNA__06310__A _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_196_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_196_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08886__A2 _02515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12458__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11979_ _05807_ _05825_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__nor2_4
X_13718_ clknet_leaf_34_clk total_design.core.data_mem.stored_read_data\[25\] net1067
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13649_ clknet_leaf_47_clk total_design.core.data_mem.data_write_adr_i\[21\] net1098
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09767__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07170_ total_design.core.regFile.register\[23\]\[12\] net681 net670 total_design.core.regFile.register\[20\]\[12\]
+ _02708_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10706__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_120_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09068__A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08023__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07377__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout317 _02287_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_4
X_09811_ net167 net2755 net440 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__mux2_1
Xfanout328 net331 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__buf_2
Xfanout339 net343 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_1
XFILLER_0_94_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11537__S net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10441__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ total_design.core.ctrl.instruction\[31\] net886 net754 total_design.core.data_cpu_o\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__a22oi_2
X_06954_ total_design.core.regFile.register\[20\]\[8\] net672 _02502_ _02504_ net688
+ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07129__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12122__A2 _05850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07316__A total_design.core.ctrl.instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09673_ _04853_ _04898_ net466 vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__mux2_1
X_06885_ _02439_ _02440_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_187_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_187_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08624_ total_design.lcd_display.cnt_20ms\[11\] total_design.lcd_display.cnt_20ms\[10\]
+ total_design.lcd_display.cnt_20ms\[13\] total_design.lcd_display.cnt_20ms\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__or4_1
XANTENNA__11881__A1 total_design.core.math.pc_val\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08555_ total_design.keypad0.key_out\[13\] net931 net932 _03861_ total_design.keypad0.key_out\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_46_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1183_A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_A _03676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07506_ total_design.core.regFile.register\[13\]\[18\] net786 net775 total_design.core.regFile.register\[22\]\[18\]
+ _03020_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__a221o_1
XANTENNA__07837__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08486_ _03817_ _03819_ _03838_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07301__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06593__C net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07437_ total_design.core.regFile.register\[25\]\[17\] net647 net624 total_design.core.regFile.register\[14\]\[17\]
+ _02950_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_21_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_99_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06890__A total_design.core.ctrl.instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07368_ _02894_ _02895_ net721 vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_165_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09107_ _04354_ _04356_ net317 vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__mux2_1
X_06319_ _01894_ _01895_ _01896_ _01897_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__nor4_1
XFILLER_0_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_111_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10616__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07299_ total_design.core.regFile.register\[16\]\[14\] _01947_ net827 total_design.core.regFile.register\[1\]\[14\]
+ _02819_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_131_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09038_ _04289_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09211__C1 _04105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold360 total_design.lcd_display.row_2\[112\] vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 total_design.lcd_display.row_2\[105\] vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 total_design.lcd_display.row_2\[70\] vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _05228_ _05233_ _05230_ _05229_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__o211ai_1
Xhold393 total_design.lcd_display.row_2\[22\] vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09706__A _03602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_X net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06576__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11447__S net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 net841 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__buf_4
Xfanout851 net852 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10351__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout862 net864 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09425__B net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout873 _01934_ vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_16
Xfanout884 _03671_ vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12113__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout895 net896 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__buf_2
XFILLER_0_172_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12951_ clknet_leaf_123_clk _00418_ net1166 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_178_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_178_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1060 total_design.core.regFile.register\[14\]\[29\] vssd1 vssd1 vccd1 vccd1 net2376
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 total_design.core.regFile.register\[26\]\[30\] vssd1 vssd1 vccd1 vccd1 net2387
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11902_ _03981_ _03983_ _05778_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__o21a_1
Xhold1082 total_design.core.regFile.register\[3\]\[21\] vssd1 vssd1 vccd1 vccd1 net2398
+ sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ clknet_leaf_138_clk _00349_ net1184 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1093 total_design.core.regFile.register\[26\]\[16\] vssd1 vssd1 vccd1 vccd1 net2409
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07540__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11833_ total_design.lcd_display.currentState\[1\] total_design.lcd_display.currentState\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_159_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14552_ net1272 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XANTENNA__07828__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11764_ net930 _01854_ _05698_ net956 net1521 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_161_Right_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09293__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13503_ clknet_leaf_181_clk _00970_ net1043 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ net195 net2552 net357 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ clknet_leaf_36_clk _01550_ net1072 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_153_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11695_ net30 net935 net878 net1792 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__o22a_1
XFILLER_0_125_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13434_ clknet_leaf_124_clk _00901_ net1187 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ net205 net2813 net476 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_102_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13365_ clknet_leaf_158_clk _00832_ net1143 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10577_ net213 net2681 net369 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12316_ _01581_ _01582_ _01580_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13296_ clknet_leaf_184_clk _00763_ net1037 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12247_ net902 _02746_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12178_ _06027_ _06028_ _06020_ _06022_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__a211oi_1
XANTENNA__11560__A0 _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ _05387_ _05376_ _05377_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__mux2_2
XANTENNA__10261__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12104__A2 _05832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_169_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_169_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_155_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06670_ net333 net332 vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__or2_1
XANTENNA__06397__D net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07531__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08340_ net1469 net938 _03704_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[27\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13194__RESET_B net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08271_ net1376 net557 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[21\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_157_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07222_ total_design.core.regFile.register\[24\]\[13\] net573 net566 total_design.core.regFile.register\[12\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07153_ _02647_ _02693_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__xor2_2
XFILLER_0_144_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10436__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11121__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07598__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07084_ total_design.core.regFile.register\[16\]\[10\] _01932_ net861 total_design.core.regFile.register\[14\]\[10\]
+ net691 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14205__Q net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1029_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06502__X _02076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout136 _05686_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout147 net148 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout489_A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout158 _05676_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_2
XANTENNA__10171__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11796__A_N net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout169 _04929_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07986_ total_design.core.regFile.register\[30\]\[28\] net839 _03480_ _03481_ _03483_
+ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09960__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07046__A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09725_ _04124_ _04943_ _04948_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__a21o_2
X_06937_ _02468_ _02488_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_87_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout656_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09656_ _04531_ _04666_ _04534_ net295 vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06868_ total_design.core.regFile.register\[18\]\[6\] net858 net844 total_design.core.regFile.register\[25\]\[6\]
+ _02424_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_26_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08607_ net1739 net342 net716 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[28\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_26_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _04463_ _04666_ _04816_ _04194_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_65_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout823_A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06730__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06799_ _02354_ _02356_ _02358_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08538_ total_design.keypad0.key_out\[13\] net932 vssd1 vssd1 vccd1 vccd1 _03887_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_102_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11015__B _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ net717 _03822_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[6\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout611_X net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10500_ net272 net2019 net483 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11480_ net1599 _05643_ net153 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__mux2_1
XANTENNA__09027__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10431_ net270 net2833 net382 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10346__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07589__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__A1 _02565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ clknet_leaf_167_clk _00617_ net1155 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10362_ net284 net2715 net484 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06797__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ total_design.lcd_display.row_1\[117\] _05814_ _05848_ total_design.lcd_display.row_2\[125\]
+ _05957_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__a221o_1
X_13081_ clknet_leaf_195_clk _00548_ net1010 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10293_ net168 net2465 net499 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__mux2_1
X_12032_ total_design.lcd_display.row_1\[114\] _05814_ _05829_ total_design.lcd_display.row_1\[106\]
+ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__a22o_1
Xhold190 net52 vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11685__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10081__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09870__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout670 net673 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11972__Y _05834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07761__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06498__C net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout681 _02038_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_8
Xfanout692 net694 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__buf_4
X_13983_ clknet_leaf_83_clk _01163_ net1241 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08994__B _03273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ clknet_leaf_200_clk _00401_ net1002 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12865_ clknet_leaf_121_clk _00332_ net1192 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11058__C1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11816_ net1844 _05709_ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__xor2_1
X_12796_ clknet_leaf_31_clk _00263_ net1060 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[23\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ net1307 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_174_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11073__A2 total_design.core.data_bus_o\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11747_ net83 net960 net293 net2785 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__a22o_1
XANTENNA__11640__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14466_ clknet_leaf_52_clk net1421 net1095 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11678_ _05643_ net1628 net131 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13417_ clknet_leaf_177_clk _00884_ net1046 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10256__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10629_ net268 net2803 net477 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__mux2_1
X_14397_ net986 total_design.keypad0.next_rows\[3\] net1085 vssd1 vssd1 vccd1 vccd1
+ net115 sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06306__Y _01885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08234__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13348_ clknet_leaf_105_clk _00815_ net1233 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13279_ clknet_leaf_183_clk _00746_ net1136 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire457_A _03131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09065__B net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ total_design.core.regFile.register\[12\]\[25\] net774 net772 total_design.core.regFile.register\[28\]\[25\]
+ _03343_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07752__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ _03273_ _03274_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09510_ _03184_ _04741_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__nor2_1
X_06722_ net551 _02263_ _02266_ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__o21a_1
XANTENNA__08249__X _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07504__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09081__A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ _04676_ _04677_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__or2_2
XFILLER_0_91_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06653_ total_design.core.regFile.register\[21\]\[2\] net597 net577 total_design.core.regFile.register\[27\]\[2\]
+ _02220_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__a221o_1
XANTENNA__06712__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09372_ _04611_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06584_ total_design.core.regFile.register\[1\]\[1\] net741 net736 net728 vssd1 vssd1
+ vccd1 vccd1 _02155_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08323_ total_design.core.data_mem.data_write_adr_reg\[19\] net546 net538 total_design.core.data_mem.data_read_adr_reg\[19\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12261__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11550__S net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout237_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08254_ net1367 net559 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[4\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_117_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07205_ _02742_ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__inv_2
XANTENNA__10166__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08185_ net891 _03512_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[28\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout404_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09955__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07136_ total_design.core.regFile.register\[4\]\[11\] net815 net776 total_design.core.regFile.register\[22\]\[11\]
+ net694 vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10961__Y _05220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11772__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07067_ total_design.core.regFile.register\[6\]\[10\] net581 _02602_ _02604_ _02611_
+ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_37_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07991__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08160__A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout773_A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07743__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout940_A _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ net749 _03467_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[27\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06951__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09708_ _03556_ _04892_ _04913_ _04931_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__o211a_1
X_10980_ _05236_ _05238_ _05212_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_104_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09639_ net507 _04866_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06703__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout826_X net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12650_ clknet_leaf_25_clk _00117_ net1106 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[28\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11601_ _05655_ net1655 net138 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__mux2_1
X_12581_ clknet_leaf_118_clk _00048_ net1169 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11460__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10263__A0 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14320_ clknet_leaf_67_clk _01481_ net1112 vssd1 vssd1 vccd1 vccd1 total_design.core.math.pc_val\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_11532_ net1600 _05670_ net147 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10802__A2 _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ clknet_leaf_106_clk _01431_ net1234 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11463_ net1532 _05663_ net155 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__mux2_1
XANTENNA__10076__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13202_ clknet_leaf_137_clk _00669_ net1180 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09865__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08759__A1 _02918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10414_ net211 net2400 net386 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14182_ clknet_leaf_79_clk net1811 net1218 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11967__Y _05829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11394_ _05602_ _05607_ _05589_ _05601_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__a211o_4
XTAP_TAPCELL_ROW_78_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13133_ clknet_leaf_6_clk _00600_ net1017 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10345_ net222 net2814 net490 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07982__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13064_ clknet_leaf_171_clk _00531_ net1056 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10276_ net228 net2467 net496 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09184__A1 _02492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12015_ total_design.lcd_display.row_2\[89\] _05837_ _05839_ total_design.lcd_display.row_1\[57\]
+ _05875_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__a221o_1
XANTENNA__13815__RESET_B net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07195__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07734__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08931__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13966_ clknet_leaf_103_clk _01146_ net1238 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07414__A _02917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12917_ clknet_leaf_159_clk _00384_ net1143 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13897_ clknet_leaf_97_clk _01077_ net1245 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08229__B net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12848_ clknet_leaf_185_clk _00315_ net1037 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10775__A total_design.core.data_bus_o\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12779_ clknet_leaf_114_clk _00246_ net1202 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12768__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14518_ net1290 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_16_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14449_ clknet_leaf_66_clk net1375 net1122 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09775__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold904 total_design.core.regFile.register\[7\]\[29\] vssd1 vssd1 vccd1 vccd1 net2220
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11102__C _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold915 total_design.core.regFile.register\[1\]\[25\] vssd1 vssd1 vccd1 vccd1 net2231
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold926 total_design.core.regFile.register\[28\]\[12\] vssd1 vssd1 vccd1 vccd1 net2242
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08899__B _02182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11754__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold937 total_design.core.regFile.register\[15\]\[30\] vssd1 vssd1 vccd1 vccd1 net2253
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 total_design.core.regFile.register\[29\]\[18\] vssd1 vssd1 vccd1 vccd1 net2264
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09990_ net281 net2546 net414 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__mux2_1
XANTENNA__10714__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold959 total_design.core.regFile.register\[11\]\[25\] vssd1 vssd1 vccd1 vccd1 net2275
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07973__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08941_ net314 _04194_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__nor2_1
X_08872_ _02112_ net462 vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__nand2_1
XANTENNA__13556__RESET_B net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07186__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07823_ _03278_ _03281_ _03326_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_84_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07754_ total_design.core.regFile.register\[29\]\[23\] net655 net592 total_design.core.regFile.register\[1\]\[23\]
+ _03260_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__a221o_1
XANTENNA__12230__A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06705_ total_design.core.regFile.register\[22\]\[3\] net674 net624 total_design.core.regFile.register\[14\]\[3\]
+ _02269_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07685_ total_design.core.regFile.register\[14\]\[22\] net862 _03193_ _03194_ vssd1
+ vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout354_A _05018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1096_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09424_ _02992_ _04659_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__xnor2_1
X_06636_ net692 _02204_ _02205_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__or3_1
XFILLER_0_149_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09355_ _02845_ net701 _04594_ net533 vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout521_A _01885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout142_X net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06567_ total_design.core.regFile.register\[20\]\[1\] _01992_ _02130_ _02133_ _02136_
+ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1263_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08306_ net1479 net940 _03687_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[10\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09286_ _04441_ _04528_ net332 vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07110__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06498_ net745 net737 net730 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11993__B1 _05840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08237_ net1420 net543 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[20\]
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_X net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09685__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08168_ _02021_ _02694_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[11\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_160_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout890_A _02022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10691__Y _05017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07119_ total_design.core.regFile.register\[10\]\[11\] net619 net570 total_design.core.regFile.register\[17\]\[11\]
+ _02660_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__a221o_1
XANTENNA__10624__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08099_ total_design.core.regFile.register\[26\]\[30\] net646 _03588_ _03591_ vssd1
+ vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10130_ net251 net2736 net400 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10061_ net266 net2587 net406 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06924__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__S net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13820_ clknet_leaf_113_clk total_design.core.data_mem.data_cpu_i\[29\] net1206 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[29\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_162_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09469__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13751_ clknet_leaf_113_clk total_design.core.data_mem.stored_write_data\[26\] net1207
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[26\] sky130_fd_sc_hd__dfrtp_1
X_10963_ _05185_ _05191_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_82_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08141__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12702_ clknet_leaf_175_clk _00169_ net1053 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13682_ clknet_leaf_47_clk total_design.core.data_mem.data_read_adr_i\[22\] net1098
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10894_ _05135_ _05139_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_156_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12633_ clknet_leaf_188_clk _00100_ net1009 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12564_ net1459 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14303_ clknet_leaf_104_clk _00017_ net1235 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11515_ net1580 _05646_ net151 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__mux2_1
X_12495_ net975 total_design.core.instr_mem.instruction_i\[11\] vssd1 vssd1 vccd1
+ vccd1 _01702_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14234_ clknet_leaf_57_clk _01414_ net1118 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12528__A2 total_design.core.ctrl.instruction\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_44_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11446_ net1716 _05648_ net158 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06207__A2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10534__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14165_ clknet_leaf_30_clk _01345_ net1060 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11377_ total_design.core.data_bus_o\[20\] net700 _05610_ vssd1 vssd1 vccd1 vccd1
+ _05636_ sky130_fd_sc_hd__a21o_2
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13116_ clknet_leaf_32_clk _00583_ net1061 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10328_ _04113_ _04118_ _05002_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__or3_1
X_14096_ clknet_leaf_110_clk _01276_ net1226 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[50\]
+ sky130_fd_sc_hd__dfrtp_1
X_13047_ clknet_leaf_164_clk _00514_ net1165 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10259_ _04929_ net2218 net500 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__mux2_1
XANTENNA__07168__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07707__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1240 net1264 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_4
Xfanout1251 net1252 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__buf_2
Xfanout1262 net1263 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06915__B1 _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13791__D total_design.core.data_mem.data_cpu_i\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11218__X _05477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13949_ clknet_leaf_92_clk _01129_ net1258 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_73_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_147_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07470_ _02949_ _02992_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_159_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07340__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06421_ net921 net916 net908 vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__and3_4
XANTENNA__10709__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10227__B1 total_design.core.instr_fetch vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09140_ _04235_ _04240_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__or2_1
X_06352_ total_design.core.ctrl.instruction\[20\] total_design.core.ctrl.instruction\[21\]
+ net951 net950 net952 vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__o221a_2
XANTENNA__09093__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_62_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06283_ total_design.core.instr_mem.instruction_adr_i\[6\] total_design.core.instr_mem.instruction_adr_stored\[6\]
+ net984 vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__mux2_1
X_09071_ _04265_ _04270_ net467 vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08022_ total_design.core.regFile.register\[23\]\[29\] net810 _03517_ vssd1 vssd1
+ vccd1 vccd1 _03518_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold701 total_design.core.regFile.register\[8\]\[26\] vssd1 vssd1 vccd1 vccd1 net2017
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold712 total_design.core.regFile.register\[24\]\[6\] vssd1 vssd1 vccd1 vccd1 net2028
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 total_design.core.regFile.register\[14\]\[17\] vssd1 vssd1 vccd1 vccd1 net2039
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09396__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold734 total_design.core.regFile.register\[13\]\[27\] vssd1 vssd1 vccd1 vccd1 net2050
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10444__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold745 total_design.core.regFile.register\[27\]\[17\] vssd1 vssd1 vccd1 vccd1 net2061
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 total_design.core.regFile.register\[6\]\[3\] vssd1 vssd1 vccd1 vccd1 net2072
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold767 total_design.core.regFile.register\[21\]\[5\] vssd1 vssd1 vccd1 vccd1 net2083
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 total_design.core.regFile.register\[26\]\[12\] vssd1 vssd1 vccd1 vccd1 net2094
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09973_ net203 net2110 net419 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__mux2_1
Xhold789 total_design.core.regFile.register\[7\]\[30\] vssd1 vssd1 vccd1 vccd1 net2105
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ _04176_ _04177_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12152__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1109_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1401 total_design.core.regFile.register\[2\]\[21\] vssd1 vssd1 vccd1 vccd1 net2717
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_71_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1412 total_design.core.regFile.register\[3\]\[14\] vssd1 vssd1 vccd1 vccd1 net2728
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08855_ _04096_ _04102_ _04109_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__a21o_1
XFILLER_0_157_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1423 total_design.core.regFile.register\[6\]\[28\] vssd1 vssd1 vccd1 vccd1 net2739
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06906__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1434 total_design.core.regFile.register\[11\]\[15\] vssd1 vssd1 vccd1 vccd1 net2750
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout569_A _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1445 total_design.core.regFile.register\[6\]\[8\] vssd1 vssd1 vccd1 vccd1 net2761
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07806_ total_design.core.regFile.register\[25\]\[24\] net648 _03309_ _03310_ net687
+ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1456 total_design.core.regFile.register\[1\]\[27\] vssd1 vssd1 vccd1 vccd1 net2772
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1467 total_design.core.regFile.register\[14\]\[19\] vssd1 vssd1 vccd1 vccd1 net2783
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08786_ _02565_ total_design.core.data_mem.data_cpu_i\[9\] _04040_ vssd1 vssd1 vccd1
+ vccd1 _04041_ sky130_fd_sc_hd__a21oi_1
Xhold1478 total_design.core.regFile.register\[16\]\[21\] vssd1 vssd1 vccd1 vccd1 net2794
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_140_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1489 total_design.core.regFile.register\[22\]\[6\] vssd1 vssd1 vccd1 vccd1 net2805
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_140_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ _03240_ _03242_ _03243_ _03244_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout736_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08123__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07989__A _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07668_ net554 total_design.core.ctrl.imm_32\[21\] vssd1 vssd1 vccd1 vccd1 _03179_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07331__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09407_ _04596_ _04644_ net460 vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__mux2_1
X_06619_ total_design.core.regFile.register\[2\]\[2\] net784 vssd1 vssd1 vccd1 vccd1
+ _02189_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10619__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06685__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07599_ total_design.core.regFile.register\[25\]\[20\] net842 net786 total_design.core.regFile.register\[13\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout903_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1266_X net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10218__A0 _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_80_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09338_ _02791_ net504 net446 _02793_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11966__B1 _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ net312 _04306_ _04191_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11300_ _05556_ _05558_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12280_ net993 _06117_ _06118_ _06119_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13876__D total_design.core.ctrl.imm_32\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11231_ _05389_ _05485_ _05489_ _05483_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__o22ai_2
XTAP_TAPCELL_ROW_75_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10354__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07937__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _05415_ _05417_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_112_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10113_ net182 net2577 net403 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_164_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11093_ _05345_ _05348_ _05349_ _05351_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__or4_1
XANTENNA__12143__B1 _05839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09444__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ net192 net2696 net411 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__mux2_1
Xhold50 total_design.core.data_mem.data_bus_i_reg\[3\] vssd1 vssd1 vccd1 vccd1 net1366
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 total_design.core.math.pc_val\[29\] vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold72 total_design.core.data_mem.data_cpu_i_reg\[10\] vssd1 vssd1 vccd1 vccd1 net1388
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 total_design.core.instr_mem.instruction_adr_stored\[2\] vssd1 vssd1 vccd1
+ vccd1 net1399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 total_design.core.instr_mem.instruction_adr_stored\[3\] vssd1 vssd1 vccd1
+ vccd1 net1410 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ clknet_leaf_76_clk total_design.core.data_mem.data_cpu_i\[12\] net1213 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[12\] sky130_fd_sc_hd__dfrtp_1
X_11995_ total_design.lcd_display.row_1\[120\] _05843_ _05847_ total_design.lcd_display.row_2\[32\]
+ _05856_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_55_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08114__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13734_ clknet_leaf_75_clk total_design.core.data_mem.stored_write_data\[9\] net1215
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[9\] sky130_fd_sc_hd__dfrtp_1
X_10946_ _05169_ _05204_ _05124_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07322__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_119_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13665_ clknet_leaf_61_clk total_design.core.data_mem.data_read_adr_i\[5\] net1129
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[5\] sky130_fd_sc_hd__dfrtp_1
X_10877_ _05111_ _05115_ _05117_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__and3_1
XANTENNA__10529__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10209__A0 _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12616_ clknet_leaf_24_clk _00083_ net1056 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13596_ clknet_leaf_62_clk net1344 net1125 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06308__A _01852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12547_ net1431 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12478_ net982 total_design.core.ctrl.instruction\[2\] net883 _01693_ vssd1 vssd1
+ vccd1 vccd1 _01541_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_3 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14217_ clknet_leaf_59_clk _01397_ net1127 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11429_ _05323_ _05354_ _05678_ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__a21boi_1
XANTENNA__10264__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08242__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07928__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14148_ clknet_leaf_43_clk _01328_ net1083 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13148__RESET_B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11884__A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06600__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14079_ clknet_leaf_83_clk _01259_ net1242 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_06970_ total_design.core.regFile.register\[1\]\[8\] net829 net812 total_design.core.regFile.register\[23\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__a22o_1
XANTENNA__12134__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1070 net1072 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__clkbuf_4
Xfanout1081 net1135 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_2
X_08640_ total_design.lcd_display.cnt_500hz\[3\] _03921_ vssd1 vssd1 vccd1 vccd1 _03929_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_174_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1092 net1096 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07561__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08571_ net1832 net339 net718 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[26\]
+ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_46_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09302__A1 _02666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07522_ total_design.core.ctrl.instruction\[19\] _02994_ vssd1 vssd1 vccd1 vccd1
+ _03041_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07453_ total_design.core.regFile.register\[5\]\[17\] net806 _02972_ vssd1 vssd1
+ vccd1 vccd1 _02977_ sky130_fd_sc_hd__a21o_1
XANTENNA__10439__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06404_ _01739_ net918 _01948_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__and3_4
XFILLER_0_88_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07384_ total_design.core.regFile.register\[29\]\[16\] net656 net634 total_design.core.regFile.register\[16\]\[16\]
+ _02910_ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09123_ net905 _04371_ _04372_ net752 _01752_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__o32a_1
X_06335_ _01910_ _01913_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10620__A0 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1059_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09529__A _03178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09054_ _04304_ _04305_ net324 vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__mux2_1
X_06266_ _01840_ _01841_ _01843_ _01844_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__o22a_1
XFILLER_0_130_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08005_ _03495_ _03497_ _03499_ _03501_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__or4_1
Xhold520 net45 vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10174__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06197_ _01762_ _01772_ _01774_ _01776_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__o22a_1
XANTENNA__13571__RESET_B net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold531 total_design.data_in_BUS\[17\] vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold542 total_design.lcd_display.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09963__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold553 total_design.core.regFile.register\[5\]\[1\] vssd1 vssd1 vccd1 vccd1 net1869
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold564 _05716_ vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 total_design.data_in_BUS\[29\] vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 total_design.core.regFile.register\[7\]\[13\] vssd1 vssd1 vccd1 vccd1 net1902
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 total_design.core.regFile.register\[4\]\[6\] vssd1 vssd1 vccd1 vccd1 net1913
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09956_ net280 total_design.core.regFile.register\[23\]\[4\] net418 vssd1 vssd1 vccd1
+ vccd1 _00267_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12125__B1 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08907_ net471 _03506_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__or2_1
X_09887_ net270 net2816 net427 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__mux2_1
Xhold1220 total_design.core.regFile.register\[11\]\[3\] vssd1 vssd1 vccd1 vccd1 net2536
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout853_A _01949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08344__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09541__A1 _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1231 total_design.core.regFile.register\[4\]\[19\] vssd1 vssd1 vccd1 vccd1 net2547
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 total_design.core.regFile.register\[24\]\[18\] vssd1 vssd1 vccd1 vccd1 net2558
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08838_ _04013_ _04092_ _04011_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1253 total_design.core.regFile.register\[21\]\[23\] vssd1 vssd1 vccd1 vccd1 net2569
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06400__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1264 total_design.core.regFile.register\[3\]\[6\] vssd1 vssd1 vccd1 vccd1 net2580
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 total_design.core.regFile.register\[3\]\[22\] vssd1 vssd1 vccd1 vccd1 net2591
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12428__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1286 total_design.core.regFile.register\[30\]\[19\] vssd1 vssd1 vccd1 vccd1 net2602
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1297 total_design.core.regFile.register\[24\]\[21\] vssd1 vssd1 vccd1 vccd1 net2613
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout641_X net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ total_design.core.data_mem.data_cpu_i\[31\] net305 vssd1 vssd1 vccd1 vccd1
+ _04024_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_37_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10800_ _01728_ _05030_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__nor2_2
XFILLER_0_135_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11780_ net1838 net953 _05694_ _01826_ vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10731_ net2570 net356 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__and2_1
XANTENNA__10349__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout906_X net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13450_ clknet_leaf_20_clk _00917_ net1050 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10662_ net268 net2294 net362 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12401_ _01658_ _01659_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13381_ clknet_leaf_118_clk _00848_ net1160 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08804__B1 total_design.core.data_mem.data_cpu_i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10593_ net286 net2117 net365 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__mux2_1
X_12332_ total_design.core.math.pc_val\[21\] total_design.core.program_count.imm_val_reg\[21\]
+ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07083__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12263_ net900 _02796_ net525 vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06830__A2 _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10084__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14002_ clknet_leaf_86_clk _01182_ net1247 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11214_ _05451_ _05461_ _05466_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__or3_2
XANTENNA__09873__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11975__Y _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12194_ total_design.core.math.pc_val\[6\] total_design.core.program_count.imm_val_reg\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__and2_1
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__clkbuf_4
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08997__B _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__clkbuf_4
X_11145_ _05402_ _05403_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__nand2_1
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12116__B1 _05838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07791__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
X_11076_ total_design.core.data_bus_o\[20\] total_design.core.data_bus_o\[28\] net695
+ _05046_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ net265 net2764 net410 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__mux2_1
XANTENNA__07543__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06897__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_127_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_28_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11978_ _05813_ _05820_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__nor2_4
X_10929_ _05185_ _05186_ _05181_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__or3b_2
XANTENNA_clkbuf_leaf_152_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06649__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13717_ clknet_leaf_27_clk total_design.core.data_mem.stored_read_data\[24\] net1077
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[24\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10259__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06309__Y _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13648_ clknet_leaf_50_clk total_design.core.data_mem.data_write_adr_i\[20\] net1102
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[20\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13579_ clknet_leaf_32_clk total_design.core.data_mem.data_bus_i\[15\] net1062 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_167_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07074__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06325__X _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06821__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12355__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09783__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09810_ net169 net2153 net438 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10722__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout318 net321 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_2
Xfanout329 net330 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__buf_2
XANTENNA__12107__B1 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ total_design.core.math.pc_val\[31\] _04944_ vssd1 vssd1 vccd1 vccd1 _04964_
+ sky130_fd_sc_hd__xnor2_2
X_06953_ total_design.core.regFile.register\[21\]\[8\] net599 net568 total_design.core.regFile.register\[12\]\[8\]
+ _02503_ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08326__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ net335 _03459_ _04161_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__o21ai_1
X_06884_ _02438_ net311 vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__nand2b_1
XANTENNA__06995__X total_design.core.ctrl.imm_32\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07534__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_145_Left_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08623_ total_design.lcd_display.cnt_20ms\[15\] total_design.lcd_display.cnt_20ms\[14\]
+ total_design.lcd_display.cnt_20ms\[17\] total_design.lcd_display.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_19_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout267_A _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ net717 _03901_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[12\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07505_ total_design.core.regFile.register\[24\]\[18\] net790 net767 total_design.core.regFile.register\[7\]\[18\]
+ _03025_ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__a221o_1
X_08485_ _03836_ _03837_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10169__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout434_A _04973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1176_A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09958__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07436_ total_design.core.regFile.register\[13\]\[17\] net666 net636 total_design.core.regFile.register\[2\]\[17\]
+ _02959_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__a221o_1
XANTENNA__06593__D net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09039__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire708 _04203_ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_73_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12043__C1 _05823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout601_A _02076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07367_ total_design.core.ctrl.instruction\[16\] _02846_ vssd1 vssd1 vccd1 vccd1
+ _02895_ sky130_fd_sc_hd__nand2_1
XANTENNA__11397__A1 total_design.core.data_bus_o\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06890__B total_design.core.ctrl.instruction\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09106_ net325 _04179_ _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__a21oi_1
X_06318_ _01782_ _01788_ _01793_ _01800_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__or4b_1
XFILLER_0_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07065__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07298_ total_design.core.regFile.register\[25\]\[14\] net842 _02830_ vssd1 vssd1
+ vccd1 vccd1 _02831_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09037_ net323 _04288_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__nor2_1
X_06249_ total_design.core.instr_mem.instruction_adr_i\[13\] total_design.core.instr_mem.instruction_adr_stored\[13\]
+ net983 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06812__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold350 total_design.lcd_display.row_1\[22\] vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 total_design.lcd_display.row_2\[16\] vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold372 total_design.lcd_display.row_2\[47\] vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold383 total_design.lcd_display.row_2\[17\] vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 total_design.lcd_display.row_2\[127\] vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10632__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout830 _01961_ vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__buf_4
Xfanout841 _01956_ vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__buf_4
Xfanout852 _01951_ vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09939_ net201 net2613 net423 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__mux2_1
Xfanout863 net864 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout856_X net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout874 _01934_ vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_4
Xfanout885 net887 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__buf_2
Xfanout896 net898 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__clkbuf_2
X_12950_ clknet_leaf_155_clk _00417_ net1137 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1050 total_design.core.regFile.register\[18\]\[5\] vssd1 vssd1 vccd1 vccd1 net2366
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11901_ _05778_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__inv_2
Xhold1061 total_design.core.regFile.register\[4\]\[20\] vssd1 vssd1 vccd1 vccd1 net2377
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 total_design.core.regFile.register\[2\]\[17\] vssd1 vssd1 vccd1 vccd1 net2388
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 total_design.core.regFile.register\[5\]\[24\] vssd1 vssd1 vccd1 vccd1 net2399
+ sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ clknet_leaf_150_clk _00348_ net1147 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06879__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1094 total_design.core.regFile.register\[23\]\[23\] vssd1 vssd1 vccd1 vccd1 net2410
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11463__S net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ total_design.lcd_display.currentState\[1\] total_design.lcd_display.currentState\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_29_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ net1271 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_56_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11763_ _01904_ _05697_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__and2_1
XANTENNA__10079__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10714_ net199 net2503 net359 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__mux2_1
XANTENNA__09868__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13502_ clknet_leaf_181_clk _00969_ net1044 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ clknet_leaf_37_clk _01549_ net1077 vssd1 vssd1 vccd1 vccd1 total_design.core.ctrl.instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_11694_ net29 net937 _05690_ net2031 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13433_ clknet_leaf_195_clk _00900_ net1010 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10645_ net211 net2326 net477 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13493__RESET_B net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07056__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13364_ clknet_leaf_144_clk _00831_ net1176 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10576_ net222 net2119 net372 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12315_ _01580_ _01581_ _01582_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__or3_1
XANTENNA__07461__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06803__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13295_ clknet_leaf_147_clk _00762_ net1152 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12246_ _06089_ total_design.core.math.pc_val\[11\] net527 vssd1 vssd1 vccd1 vccd1
+ _01481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11638__S net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ total_design.core.math.pc_val\[4\] total_design.core.program_count.imm_val_reg\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__or2_1
XANTENNA__09616__B _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10542__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07764__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ _05371_ _05376_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__nand2_1
XANTENNA__08308__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09505__A1 total_design.core.ctrl.instruction\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11059_ total_design.core.data_bus_o\[18\] net695 _05298_ net517 vssd1 vssd1 vccd1
+ vccd1 _05318_ sky130_fd_sc_hd__a211o_1
XANTENNA__10778__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09778__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08270_ net1392 net558 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[20\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11105__C net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06991__A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07295__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07221_ total_design.core.regFile.register\[9\]\[13\] net663 net644 total_design.core.regFile.register\[26\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10717__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07152_ _02689_ _02690_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__nand2b_2
XANTENNA__12040__A2 _05840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06341__A_N total_design.core.ctrl.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07083_ total_design.core.regFile.register\[28\]\[10\] net853 net810 total_design.core.regFile.register\[23\]\[10\]
+ _02627_ vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11548__S net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10452__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09526__B _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14369__RESET_B net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11551__A1 _05651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07755__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 net138 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_4
Xfanout148 _05683_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_4
Xfanout159 _05676_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_4
X_07985_ total_design.core.regFile.register\[19\]\[28\] net824 net791 total_design.core.regFile.register\[24\]\[28\]
+ _03482_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__a221o_1
X_09724_ total_design.core.ctrl.instruction\[30\] net889 net755 total_design.core.data_cpu_o\[30\]
+ _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__a221o_1
X_06936_ _02468_ _02488_ vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__nand2_1
XANTENNA__12500__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09655_ _04880_ _04881_ _04193_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06867_ total_design.core.regFile.register\[26\]\[6\] net871 net799 total_design.core.regFile.register\[29\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout551_A _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ net1635 net342 net716 vssd1 vssd1 vccd1 vccd1 total_design.core.data_out_INSTR\[27\]
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout649_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_26_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09586_ _04646_ _04815_ net318 vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08158__A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06798_ total_design.core.regFile.register\[19\]\[5\] net642 net590 total_design.core.regFile.register\[1\]\[5\]
+ _02357_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_65_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _03862_ _03885_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1081_X net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1499_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10200__B net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout816_A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08468_ total_design.data_in_BUS\[6\] _01888_ _03821_ net519 vssd1 vssd1 vccd1 vccd1
+ _03822_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_61_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07286__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07419_ net750 _02944_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[16\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08399_ total_design.keypad0.key_out\[13\] _03754_ vssd1 vssd1 vccd1 vccd1 _03755_
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout604_X net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10627__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10430_ net276 net2256 net382 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12031__A2 _05812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06406__A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08786__A2 total_design.core.data_mem.data_cpu_i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10361_ _04971_ _04972_ _05002_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__or3_4
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12100_ total_design.lcd_display.row_2\[77\] _05806_ _05837_ total_design.lcd_display.row_2\[93\]
+ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__a22o_1
XANTENNA__07994__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11790__B2 _01793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13080_ clknet_leaf_136_clk _00547_ net1179 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10292_ net170 net2376 net496 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__mux2_1
XANTENNA__11781__A2_N _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout973_X net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11458__S net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ total_design.lcd_display.row_1\[90\] _05812_ _05841_ total_design.lcd_display.row_1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold180 total_design.core.data_mem.data_cpu_i_reg\[28\] vssd1 vssd1 vccd1 vccd1 net1496
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10362__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold191 net110 vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11542__A1 _05609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout660 net662 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06954__D1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout671 net673 vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_4
XANTENNA__12098__A2 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout682 _02035_ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_16
X_13982_ clknet_leaf_100_clk _01162_ net1254 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout693 net694 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ clknet_leaf_117_clk _00400_ net1160 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12864_ clknet_leaf_201_clk _00331_ net1003 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11815_ _05709_ _05710_ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__nor2_1
X_12795_ clknet_leaf_144_clk _00262_ net1174 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13674__RESET_B net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11746_ net1669 net958 net290 total_design.core.data_bus_o\[18\] vssd1 vssd1 vccd1
+ vccd1 _01374_ sky130_fd_sc_hd__a22o_1
X_14534_ net1306 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XFILLER_0_138_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07277__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11073__A3 total_design.core.data_bus_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14465_ clknet_leaf_52_clk net1423 net1095 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11677_ _05648_ net1779 net132 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10537__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10628_ net278 net2079 net477 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13416_ clknet_leaf_171_clk _00883_ net1057 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07029__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14396_ net986 total_design.keypad0.next_rows\[2\] net1085 vssd1 vssd1 vccd1 vccd1
+ net114 sky130_fd_sc_hd__dfstp_1
XANTENNA__12022__A2 _05819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13347_ clknet_leaf_5_clk _00814_ net1024 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10559_ _04984_ net532 vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__nand2_4
XFILLER_0_11_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07985__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09627__A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11876__B net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13278_ clknet_leaf_175_clk _00745_ net1052 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12229_ total_design.core.math.pc_val\[9\] net527 _06074_ vssd1 vssd1 vccd1 vccd1
+ _01479_ sky130_fd_sc_hd__a21o_1
XANTENNA__10272__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07418__Y _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11533__A1 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07770_ _03274_ _03273_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__and2b_1
XANTENNA__12089__A2 _05810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06721_ total_design.core.regFile.register\[0\]\[3\] net684 _02280_ _02285_ vssd1
+ vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__o22a_4
XANTENNA__09362__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ total_design.core.math.pc_val\[17\] _04651_ vssd1 vssd1 vccd1 vccd1 _04677_
+ sky130_fd_sc_hd__nor2_1
X_06652_ total_design.core.regFile.register\[19\]\[2\] net640 net592 total_design.core.regFile.register\[1\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09371_ _04609_ _04610_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_82_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06583_ total_design.core.regFile.register\[24\]\[1\] net746 net739 net723 vssd1
+ vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__and4_1
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08322_ net1458 net939 _03695_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_data_adr\[18\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07268__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09301__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08253_ net1359 net559 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_write_data\[3\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__10447__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07204_ _02740_ _02741_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__nor2_4
XFILLER_0_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08184_ net890 _03467_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[27\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__12013__A2 _05835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06228__B1 net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07135_ total_design.core.regFile.register\[8\]\[11\] net802 _02676_ vssd1 vssd1
+ vccd1 vccd1 _02677_ sky130_fd_sc_hd__a21o_1
XFILLER_0_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1041_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1139_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07066_ _02606_ _02608_ _02610_ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__or3_1
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07440__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10182__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08160__B _02292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11524__A1 _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07728__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09971__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout766_A _01997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _03465_ _03466_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_96_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06919_ total_design.core.regFile.register\[9\]\[7\] _01951_ net841 total_design.core.regFile.register\[30\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__a22o_1
X_09707_ net306 _03552_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__nand2b_1
X_07899_ total_design.core.regFile.register\[9\]\[26\] net664 net621 total_design.core.regFile.register\[4\]\[26\]
+ _03398_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09638_ total_design.core.data_cpu_o\[26\] net756 _04860_ _04865_ vssd1 vssd1 vccd1
+ vccd1 _04866_ sky130_fd_sc_hd__a211o_4
XANTENNA__07900__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09569_ total_design.core.math.pc_val\[23\] _04777_ vssd1 vssd1 vccd1 vccd1 _04800_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout819_X net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ _05679_ net1629 net139 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12580_ clknet_leaf_106_clk _00047_ net1223 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13879__D total_design.core.ctrl.imm_32\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11531_ net1517 _05667_ net145 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__mux2_1
XANTENNA__10357__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14250_ clknet_leaf_106_clk _01430_ net1234 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11462_ net1527 _05627_ net154 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12004__A2 _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13201_ clknet_leaf_150_clk _00668_ net1147 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10413_ net218 net2129 net388 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__mux2_1
XANTENNA__08759__A2 total_design.core.data_mem.data_cpu_i\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14181_ clknet_leaf_79_clk net1754 net1218 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
X_11393_ _05575_ net510 _05036_ _05608_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13132_ clknet_leaf_165_clk _00599_ net1158 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10344_ net226 net2850 net490 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__mux2_1
XANTENNA__07431__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10092__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13063_ clknet_leaf_174_clk _00530_ net1054 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10275_ net238 net2337 net498 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__mux2_1
XANTENNA__11515__A1 _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ total_design.lcd_display.row_1\[105\] _05829_ _05840_ total_design.lcd_display.row_1\[49\]
+ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__a22o_1
XANTENNA__09881__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09184__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11983__Y _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08931__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout490 net491 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_8
X_13965_ clknet_leaf_91_clk _01145_ net1262 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_12916_ clknet_leaf_144_clk _00383_ net1176 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[20\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07498__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13896_ clknet_leaf_74_clk _01076_ net1220 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ clknet_leaf_147_clk _00314_ net1177 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[22\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11651__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12778_ clknet_leaf_25_clk _00245_ net1106 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[24\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14517_ net1289 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08998__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10267__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11729_ net84 net960 net293 net2704 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08245__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14448_ clknet_leaf_66_clk net1411 net1122 vssd1 vssd1 vccd1 vccd1 total_design.core.instr_mem.instruction_adr_i\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10791__A total_design.core.data_bus_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14379_ clknet_leaf_187_clk _01520_ net1029 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[31\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold905 total_design.core.regFile.register\[26\]\[8\] vssd1 vssd1 vccd1 vccd1 net2221
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07958__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold916 total_design.core.regFile.register\[9\]\[7\] vssd1 vssd1 vccd1 vccd1 net2232
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__A1 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold927 total_design.core.regFile.register\[25\]\[27\] vssd1 vssd1 vccd1 vccd1 net2243
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__B2 total_design.core.data_bus_o\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold938 total_design.core.regFile.register\[8\]\[9\] vssd1 vssd1 vccd1 vccd1 net2254
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold949 total_design.core.regFile.register\[8\]\[13\] vssd1 vssd1 vccd1 vccd1 net2265
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06630__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08940_ _02338_ _04104_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__or2_4
XANTENNA__11506__A1 _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09791__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09175__A2 _04414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08871_ net967 _04123_ _01921_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__o21ai_1
X_07822_ _03278_ _03281_ _03326_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_32_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07753_ total_design.core.regFile.register\[7\]\[23\] net651 net569 total_design.core.regFile.register\[17\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08135__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06704_ total_design.core.regFile.register\[5\]\[3\] net628 net585 total_design.core.regFile.register\[28\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07489__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07684_ total_design.core.regFile.register\[30\]\[22\] net839 net787 total_design.core.regFile.register\[13\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__a22o_1
XANTENNA__12482__A2 total_design.core.ctrl.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09423_ _02992_ _04658_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__and2_1
X_06635_ total_design.core.regFile.register\[12\]\[2\] net774 net772 total_design.core.regFile.register\[28\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11561__S net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1089_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ _04592_ _04593_ net701 vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__a21oi_1
X_06566_ total_design.core.regFile.register\[6\]\[1\] net764 _02131_ _02132_ _02134_
+ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__a2111o_1
X_08305_ total_design.core.data_mem.data_write_adr_reg\[10\] net548 net540 total_design.core.data_mem.data_read_adr_reg\[10\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10177__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ _04527_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06497_ total_design.core.regFile.register\[11\]\[0\] net740 net732 net723 vssd1
+ vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout514_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout135_X net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09966__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08236_ net1436 net543 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[19\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_145_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07661__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08167_ net892 _02640_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_i\[10\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07949__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11745__B2 total_design.core.data_bus_o\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ total_design.core.regFile.register\[19\]\[11\] net643 net627 total_design.core.regFile.register\[14\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08171__A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08098_ total_design.core.regFile.register\[14\]\[30\] net626 _03589_ _03590_ vssd1
+ vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__a211o_1
XANTENNA__06621__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07049_ total_design.core.regFile.register\[5\]\[10\] net628 net601 total_design.core.regFile.register\[31\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1211_X net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ net272 net2123 net408 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08913__A2 _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10640__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09206__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10962_ net521 _05220_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__nand2_2
X_13750_ clknet_leaf_72_clk total_design.core.data_mem.stored_write_data\[25\] net1205
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11681__A0 _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06688__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12701_ clknet_leaf_10_clk _00168_ net1019 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[26\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07885__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13681_ clknet_leaf_47_clk total_design.core.data_mem.data_read_adr_i\[21\] net1098
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[21\] sky130_fd_sc_hd__dfrtp_1
X_10893_ _05129_ _05135_ _05137_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__and3_1
XANTENNA__11471__S net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14562__1282 vssd1 vssd1 vccd1 vccd1 _14562__1282/HI net1282 sky130_fd_sc_hd__conb_1
X_12632_ clknet_leaf_133_clk _00099_ net1195 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06418__X _01994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12563_ net1438 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10087__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08065__B _03559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ net1771 _05645_ net149 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__mux2_1
XANTENNA__09876__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14302_ clknet_leaf_104_clk _00016_ net1235 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11978__Y _05840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12494_ net977 total_design.core.ctrl.instruction\[10\] net882 _01701_ vssd1 vssd1
+ vccd1 vccd1 _01549_ sky130_fd_sc_hd__a22o_1
XANTENNA__07652__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14233_ clknet_leaf_57_clk _01413_ net1119 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dfrtp_1
X_11445_ net1658 _05628_ net160 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11736__B2 total_design.core.data_bus_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14164_ clknet_leaf_31_clk _01344_ net1061 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11376_ _05356_ _05462_ _05468_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__o21ai_4
XANTENNA__07404__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13695__Q total_design.core.data_cpu_o\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ net163 net2304 net493 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ clknet_leaf_143_clk _00582_ net1173 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14095_ clknet_leaf_84_clk _01275_ net1246 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06313__B _01847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13046_ clknet_leaf_156_clk _00513_ net1140 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10258_ net174 net2136 net502 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__mux2_1
Xfanout1230 net1231 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11646__S net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1241 net1243 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10550__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1252 net1264 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__clkbuf_2
X_10189_ _04280_ net2037 net390 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__mux2_1
Xfanout1263 net1264 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13948_ clknet_leaf_98_clk _01128_ net1242 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09865__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11672__A0 _05652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06679__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10786__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13879_ clknet_leaf_26_clk total_design.core.ctrl.imm_32\[18\] net1080 vssd1 vssd1
+ vccd1 vccd1 total_design.core.program_count.imm_val_reg\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06420_ net923 net912 net908 vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10227__A1 total_design.core.ctrl.instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07628__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06351_ _01736_ _01737_ _01917_ _01920_ _01915_ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09786__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09070_ net467 _04262_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__nand2_1
X_06282_ total_design.core.data_adr_o\[4\] _01860_ net964 vssd1 vssd1 vccd1 vccd1
+ _01861_ sky130_fd_sc_hd__mux2_2
XANTENNA__07643__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08021_ total_design.core.regFile.register\[26\]\[29\] net869 net786 total_design.core.regFile.register\[13\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06851__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11410__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold702 total_design.core.regFile.register\[10\]\[2\] vssd1 vssd1 vccd1 vccd1 net2018
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold713 total_design.core.regFile.register\[23\]\[12\] vssd1 vssd1 vccd1 vccd1 net2029
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08053__C1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1__f_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold724 total_design.core.regFile.register\[11\]\[9\] vssd1 vssd1 vccd1 vccd1 net2040
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 total_design.core.regFile.register\[5\]\[30\] vssd1 vssd1 vccd1 vccd1 net2051
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 total_design.core.regFile.register\[23\]\[15\] vssd1 vssd1 vccd1 vccd1 net2062
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 total_design.core.regFile.register\[10\]\[29\] vssd1 vssd1 vccd1 vccd1 net2073
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 total_design.core.regFile.register\[17\]\[6\] vssd1 vssd1 vccd1 vccd1 net2084
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09972_ net208 net2800 net418 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__mux2_1
Xhold779 total_design.core.regFile.register\[26\]\[28\] vssd1 vssd1 vccd1 vccd1 net2095
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08923_ net473 net299 vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11556__S net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1402 total_design.keypad0.key_counter\[2\] vssd1 vssd1 vccd1 vccd1 net2718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1413 total_design.core.regFile.register\[19\]\[6\] vssd1 vssd1 vccd1 vccd1 net2729
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08854_ _04096_ _04099_ _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout1004_A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1424 total_design.core.regFile.register\[22\]\[13\] vssd1 vssd1 vccd1 vccd1 net2740
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1435 total_design.core.regFile.register\[25\]\[24\] vssd1 vssd1 vccd1 vccd1 net2751
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1446 total_design.core.regFile.register\[26\]\[10\] vssd1 vssd1 vccd1 vccd1 net2762
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07805_ total_design.core.regFile.register\[23\]\[24\] net679 net617 total_design.core.regFile.register\[10\]\[24\]
+ _03304_ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08785_ _02515_ total_design.core.data_mem.data_cpu_i\[8\] vssd1 vssd1 vccd1 vccd1
+ _04040_ sky130_fd_sc_hd__and2b_1
Xhold1457 total_design.core.regFile.register\[4\]\[14\] vssd1 vssd1 vccd1 vccd1 net2773
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1468 total_design.core.regFile.register\[6\]\[23\] vssd1 vssd1 vccd1 vccd1 net2784
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1479 total_design.core.regFile.register\[16\]\[13\] vssd1 vssd1 vccd1 vccd1 net2795
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout464_A _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07736_ total_design.core.regFile.register\[18\]\[23\] net860 net830 total_design.core.regFile.register\[1\]\[23\]
+ _03235_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__a221o_1
XANTENNA__06596__D net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11663__A0 _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ net299 vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout631_A _02062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06618_ net751 _02188_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[1\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09406_ net337 _02918_ _04130_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08166__A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09608__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07598_ total_design.core.regFile.register\[0\]\[20\] net682 _03108_ _03111_ vssd1
+ vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__o22a_4
XANTENNA__07882__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06549_ total_design.core.regFile.register\[9\]\[1\] net920 net913 net909 vssd1 vssd1
+ vccd1 vccd1 _02122_ sky130_fd_sc_hd__and4_1
X_09337_ net314 _04384_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09268_ _02634_ net446 _04509_ _04511_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__o211a_1
XANTENNA__07634__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08219_ net1353 net545 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.stored_read_data\[2\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10635__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09199_ _04159_ _04434_ _04437_ net295 vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__o22a_1
XFILLER_0_50_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11230_ _05485_ _05486_ _05389_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06414__A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11161_ _05409_ _05410_ _05412_ _05418_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_112_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10112_ net185 net2036 net403 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ net352 _05095_ _05314_ _05350_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_164_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11466__S net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ net193 net2569 net410 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__mux2_1
XANTENNA__10370__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09444__B _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 total_design.core.data_mem.data_bus_i_reg\[7\] vssd1 vssd1 vccd1 vccd1 net1356
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 total_design.core.data_mem.data_cpu_i_reg\[4\] vssd1 vssd1 vccd1 vccd1 net1367
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 total_design.core.data_mem.data_bus_i_reg\[22\] vssd1 vssd1 vccd1 vccd1 net1378
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 total_design.core.math.pc_val\[30\] vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold84 total_design.core.data_mem.data_bus_i_reg\[8\] vssd1 vssd1 vccd1 vccd1 net1400
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 total_design.core.math.pc_val\[9\] vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ clknet_leaf_76_clk total_design.core.data_mem.data_cpu_i\[11\] net1214 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_cpu_i_reg\[11\] sky130_fd_sc_hd__dfrtp_1
X_11994_ total_design.lcd_display.row_2\[16\] _05845_ _05852_ total_design.lcd_display.row_2\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_4_12__f_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13733_ clknet_leaf_75_clk total_design.core.data_mem.stored_write_data\[8\] net1215
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_bus_o\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10945_ _05150_ _05175_ _05203_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06295__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13664_ clknet_leaf_61_clk total_design.core.data_mem.data_read_adr_i\[4\] net1130
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_reg\[4\] sky130_fd_sc_hd__dfrtp_1
X_10876_ _05134_ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12615_ clknet_leaf_23_clk _00082_ net1055 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13595_ clknet_leaf_27_clk total_design.core.data_mem.data_bus_i\[31\] net1076 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12546_ net1398 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10545__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12477_ net982 total_design.core.instr_mem.instruction_i\[2\] vssd1 vssd1 vccd1 vccd1
+ _01693_ sky130_fd_sc_hd__and2b_1
XANTENNA_4 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ clknet_leaf_59_clk _01396_ net1127 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfrtp_1
X_11428_ _01855_ _05024_ _05027_ _05353_ total_design.lcd_display.row_1\[105\] vssd1
+ vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__a41o_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11359_ _05440_ _05459_ _05615_ _05617_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__o2bb2ai_4
X_14147_ clknet_leaf_43_clk _01327_ net1083 vssd1 vssd1 vccd1 vccd1 total_design.data_in_BUS\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08050__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11884__B _02188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14078_ clknet_leaf_101_clk _01258_ net1237 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_2\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06611__X _02182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10280__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13029_ clknet_leaf_116_clk _00496_ net1212 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1060 net1065 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07155__A _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1071 net1072 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07010__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1083 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_4
Xfanout1093 net1096 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__buf_2
X_08570_ net2884 net339 net718 vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i\[25\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07521_ net749 _03040_ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_read_adr_i\[18\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11645__A0 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11405__A _05077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07452_ total_design.core.regFile.register\[15\]\[17\] net846 _01980_ total_design.core.regFile.register\[12\]\[17\]
+ _02971_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07864__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06403_ total_design.core.regFile.register\[11\]\[0\] net922 net915 net912 vssd1
+ vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__and4_1
XFILLER_0_57_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07383_ total_design.core.regFile.register\[7\]\[16\] net653 net605 total_design.core.regFile.register\[15\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09122_ total_design.core.math.pc_val\[4\] _04345_ vssd1 vssd1 vccd1 vccd1 _04372_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_44_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06334_ net1 _01912_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__nand2_1
XANTENNA__07077__B1 _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12070__B1 _05912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11411__Y _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06824__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09053_ _04134_ _04138_ net459 vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06265_ total_design.core.data_adr_o\[23\] net962 vssd1 vssd1 vccd1 vccd1 _01844_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10455__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11586__D_N _05675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08004_ total_design.core.regFile.register\[13\]\[28\] net667 net598 total_design.core.regFile.register\[21\]\[28\]
+ _03500_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold510 net64 vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06196_ total_design.core.mem_ctrl.state\[1\] _01725_ _01773_ vssd1 vssd1 vccd1 vccd1
+ _01776_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold521 total_design.core.regFile.register\[14\]\[1\] vssd1 vssd1 vccd1 vccd1 net1837
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 total_design.lcd_display.row_2\[108\] vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold543 _05712_ vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 total_design.lcd_display.cnt_20ms\[13\] vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08041__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold565 total_design.lcd_display.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1121_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 total_design.lcd_display.row_2\[67\] vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1219_A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold587 total_design.core.regFile.register\[1\]\[1\] vssd1 vssd1 vccd1 vccd1 net1903
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 total_design.core.regFile.register\[13\]\[25\] vssd1 vssd1 vccd1 vccd1 net1914
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14561__1281 vssd1 vssd1 vccd1 vccd1 _14561__1281/HI net1281 sky130_fd_sc_hd__conb_1
X_09955_ net270 net2042 net419 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout581_A _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout679_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10190__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ net471 net306 vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__nand2_1
X_09886_ net279 net2654 net427 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__mux2_1
Xhold1210 total_design.data_in_BUS\[2\] vssd1 vssd1 vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 total_design.core.regFile.register\[23\]\[7\] vssd1 vssd1 vccd1 vccd1 net2537
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 total_design.core.regFile.register\[14\]\[9\] vssd1 vssd1 vccd1 vccd1 net2548
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ _04004_ _04091_ _04001_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__o21ai_1
Xhold1243 total_design.core.regFile.register\[31\]\[15\] vssd1 vssd1 vccd1 vccd1 net2559
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1254 total_design.core.regFile.register\[0\]\[6\] vssd1 vssd1 vccd1 vccd1 net2570
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout846_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06400__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1265 total_design.core.regFile.register\[12\]\[14\] vssd1 vssd1 vccd1 vccd1 net2581
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1276 total_design.core.regFile.register\[28\]\[20\] vssd1 vssd1 vccd1 vccd1 net2592
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 total_design.core.regFile.register\[19\]\[31\] vssd1 vssd1 vccd1 vccd1 net2603
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12428__A2 _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1298 total_design.core.regFile.register\[28\]\[18\] vssd1 vssd1 vccd1 vccd1 net2614
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08768_ total_design.core.data_mem.data_cpu_i\[30\] _03595_ vssd1 vssd1 vccd1 vccd1
+ _04023_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11636__A0 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07719_ _03207_ _03226_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08699_ total_design.keypad0.counter\[8\] _03953_ net2480 vssd1 vssd1 vccd1 vccd1
+ _03967_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10730_ total_design.core.regFile.register\[0\]\[5\] net356 vssd1 vssd1 vccd1 vccd1
+ _01004_ sky130_fd_sc_hd__and2_1
XANTENNA__07855__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10661_ net277 net1915 net362 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12400_ _01648_ _01649_ _01650_ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07068__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12061__B1 _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13380_ clknet_leaf_130_clk _00847_ net1198 vssd1 vssd1 vccd1 vccd1 total_design.core.regFile.register\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07607__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10592_ _04986_ _05001_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__nand2_1
XANTENNA__08804__A1 total_design.core.data_mem.data_cpu_i\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08804__B2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12331_ total_design.core.math.pc_val\[21\] total_design.core.program_count.imm_val_reg\[21\]
+ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10365__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12262_ net993 _06101_ _06102_ _06103_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06144__A total_design.core.data_bus_o\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11213_ _05461_ _05466_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__nor2_1
X_14001_ clknet_leaf_94_clk _01181_ net1255 vssd1 vssd1 vccd1 vccd1 total_design.lcd_display.row_1\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12193_ total_design.core.math.pc_val\[5\] net526 _06035_ _06042_ vssd1 vssd1 vccd1
+ vccd1 _01475_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08032__A2 _01932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__clkbuf_4
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__clkbuf_4
X_11144_ _05395_ _05397_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07240__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__clkbuf_4
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__clkbuf_4
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__clkbuf_4
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11075_ net518 _05049_ _05111_ _05332_ _05333_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__o2111a_1
XANTENNA__11991__Y _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10026_ net273 net2774 net412 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11627__A0 _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08099__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11977_ _05803_ _05813_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__nor2_4
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13716_ clknet_leaf_32_clk total_design.core.data_mem.stored_read_data\[23\] net1063
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_cpu_o\[23\] sky130_fd_sc_hd__dfrtp_1
X_10928_ _05160_ _05155_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07846__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13647_ clknet_leaf_49_clk total_design.core.data_mem.data_write_adr_i\[19\] net1101
+ vssd1 vssd1 vccd1 vccd1 total_design.core.data_mem.data_write_adr_reg\[19\] sky130_fd_sc_hd__dfrtp_1
X_10859_ _05115_ _05117_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07059__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11879__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13578_ clknet_leaf_32_clk total_design.core.data_mem.data_bus_i\[14\] net1061 vssd1
+ vssd1 vccd1 vccd1 total_design.core.data_mem.data_bus_i_reg\[14\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13797__D total_design.core.data_mem.data_cpu_i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12529_ net979 total_design.core.instr_mem.instruction_i\[28\] vssd1 vssd1 vccd1
+ vccd1 _01719_ sky130_fd_sc_hd__and2b_1
XANTENNA__10275__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08253__B net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10366__A0 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout319 net321 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_4
X_06952_ total_design.core.regFile.register\[24\]\[8\] net575 net572 total_design.core.regFile.register\[17\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__a22o_1
X_09740_ _04954_ _04961_ _04962_ net450 vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__a31o_1
.ends

