module sequence_counter(
    input update_t mode,
    input logic enable,
    output logic [5:0] cmd_index;
);


endmodule