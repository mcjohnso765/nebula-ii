VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO team_03
  CLASS BLOCK ;
  FOREIGN team_03 ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 300.000 ;
  PIN ACK_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 90.250 296.000 90.530 300.000 ;
    END
  END ACK_I
  PIN ADR_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 357.510 296.000 357.790 300.000 ;
    END
  END ADR_O[0]
  PIN ADR_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 557.150 296.000 557.430 300.000 ;
    END
  END ADR_O[10]
  PIN ADR_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 537.830 296.000 538.110 300.000 ;
    END
  END ADR_O[11]
  PIN ADR_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 534.610 296.000 534.890 300.000 ;
    END
  END ADR_O[12]
  PIN ADR_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 524.950 296.000 525.230 300.000 ;
    END
  END ADR_O[13]
  PIN ADR_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 502.410 296.000 502.690 300.000 ;
    END
  END ADR_O[14]
  PIN ADR_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 473.430 296.000 473.710 300.000 ;
    END
  END ADR_O[15]
  PIN ADR_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 489.530 296.000 489.810 300.000 ;
    END
  END ADR_O[16]
  PIN ADR_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 479.870 296.000 480.150 300.000 ;
    END
  END ADR_O[17]
  PIN ADR_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 450.890 296.000 451.170 300.000 ;
    END
  END ADR_O[18]
  PIN ADR_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 457.330 296.000 457.610 300.000 ;
    END
  END ADR_O[19]
  PIN ADR_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 190.070 296.000 190.350 300.000 ;
    END
  END ADR_O[1]
  PIN ADR_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 454.110 296.000 454.390 300.000 ;
    END
  END ADR_O[20]
  PIN ADR_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 441.230 296.000 441.510 300.000 ;
    END
  END ADR_O[21]
  PIN ADR_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 421.910 296.000 422.190 300.000 ;
    END
  END ADR_O[22]
  PIN ADR_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 425.130 296.000 425.410 300.000 ;
    END
  END ADR_O[23]
  PIN ADR_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 399.370 296.000 399.650 300.000 ;
    END
  END ADR_O[24]
  PIN ADR_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 396.150 296.000 396.430 300.000 ;
    END
  END ADR_O[25]
  PIN ADR_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 383.270 296.000 383.550 300.000 ;
    END
  END ADR_O[26]
  PIN ADR_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 373.610 296.000 373.890 300.000 ;
    END
  END ADR_O[27]
  PIN ADR_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 254.470 296.000 254.750 300.000 ;
    END
  END ADR_O[28]
  PIN ADR_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 251.250 296.000 251.530 300.000 ;
    END
  END ADR_O[29]
  PIN ADR_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 595.790 296.000 596.070 300.000 ;
    END
  END ADR_O[2]
  PIN ADR_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 296.000 116.290 300.000 ;
    END
  END ADR_O[30]
  PIN ADR_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 296.000 96.970 300.000 ;
    END
  END ADR_O[31]
  PIN ADR_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 615.110 296.000 615.390 300.000 ;
    END
  END ADR_O[3]
  PIN ADR_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 618.330 296.000 618.610 300.000 ;
    END
  END ADR_O[4]
  PIN ADR_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 611.890 296.000 612.170 300.000 ;
    END
  END ADR_O[5]
  PIN ADR_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 592.570 296.000 592.850 300.000 ;
    END
  END ADR_O[6]
  PIN ADR_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 576.470 296.000 576.750 300.000 ;
    END
  END ADR_O[7]
  PIN ADR_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 573.250 296.000 573.530 300.000 ;
    END
  END ADR_O[8]
  PIN ADR_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 563.590 296.000 563.870 300.000 ;
    END
  END ADR_O[9]
  PIN CYC_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 148.210 296.000 148.490 300.000 ;
    END
  END CYC_O
  PIN DAT_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END DAT_I[0]
  PIN DAT_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END DAT_I[10]
  PIN DAT_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END DAT_I[11]
  PIN DAT_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END DAT_I[12]
  PIN DAT_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END DAT_I[13]
  PIN DAT_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END DAT_I[14]
  PIN DAT_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END DAT_I[15]
  PIN DAT_I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END DAT_I[16]
  PIN DAT_I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END DAT_I[17]
  PIN DAT_I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END DAT_I[18]
  PIN DAT_I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END DAT_I[19]
  PIN DAT_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END DAT_I[1]
  PIN DAT_I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END DAT_I[20]
  PIN DAT_I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END DAT_I[21]
  PIN DAT_I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END DAT_I[22]
  PIN DAT_I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END DAT_I[23]
  PIN DAT_I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END DAT_I[24]
  PIN DAT_I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END DAT_I[25]
  PIN DAT_I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END DAT_I[26]
  PIN DAT_I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END DAT_I[27]
  PIN DAT_I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END DAT_I[28]
  PIN DAT_I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END DAT_I[29]
  PIN DAT_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END DAT_I[2]
  PIN DAT_I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END DAT_I[30]
  PIN DAT_I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END DAT_I[31]
  PIN DAT_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END DAT_I[3]
  PIN DAT_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END DAT_I[4]
  PIN DAT_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END DAT_I[5]
  PIN DAT_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END DAT_I[6]
  PIN DAT_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END DAT_I[7]
  PIN DAT_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END DAT_I[8]
  PIN DAT_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END DAT_I[9]
  PIN DAT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 431.570 296.000 431.850 300.000 ;
    END
  END DAT_O[0]
  PIN DAT_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 244.810 296.000 245.090 300.000 ;
    END
  END DAT_O[10]
  PIN DAT_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 151.430 296.000 151.710 300.000 ;
    END
  END DAT_O[11]
  PIN DAT_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 183.630 296.000 183.910 300.000 ;
    END
  END DAT_O[12]
  PIN DAT_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 512.070 296.000 512.350 300.000 ;
    END
  END DAT_O[13]
  PIN DAT_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 541.050 296.000 541.330 300.000 ;
    END
  END DAT_O[14]
  PIN DAT_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 689.170 296.000 689.450 300.000 ;
    END
  END DAT_O[15]
  PIN DAT_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 666.630 296.000 666.910 300.000 ;
    END
  END DAT_O[16]
  PIN DAT_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 579.690 296.000 579.970 300.000 ;
    END
  END DAT_O[17]
  PIN DAT_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 692.390 296.000 692.670 300.000 ;
    END
  END DAT_O[18]
  PIN DAT_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 389.710 296.000 389.990 300.000 ;
    END
  END DAT_O[19]
  PIN DAT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 296.000 113.070 300.000 ;
    END
  END DAT_O[1]
  PIN DAT_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 685.950 296.000 686.230 300.000 ;
    END
  END DAT_O[20]
  PIN DAT_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 695.610 296.000 695.890 300.000 ;
    END
  END DAT_O[21]
  PIN DAT_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 560.370 296.000 560.650 300.000 ;
    END
  END DAT_O[22]
  PIN DAT_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 296.000 145.270 300.000 ;
    END
  END DAT_O[23]
  PIN DAT_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 222.270 296.000 222.550 300.000 ;
    END
  END DAT_O[24]
  PIN DAT_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 212.610 296.000 212.890 300.000 ;
    END
  END DAT_O[25]
  PIN DAT_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 405.810 296.000 406.090 300.000 ;
    END
  END DAT_O[26]
  PIN DAT_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 141.770 296.000 142.050 300.000 ;
    END
  END DAT_O[27]
  PIN DAT_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 196.510 296.000 196.790 300.000 ;
    END
  END DAT_O[28]
  PIN DAT_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 180.410 296.000 180.690 300.000 ;
    END
  END DAT_O[29]
  PIN DAT_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 669.850 296.000 670.130 300.000 ;
    END
  END DAT_O[2]
  PIN DAT_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 167.530 296.000 167.810 300.000 ;
    END
  END DAT_O[30]
  PIN DAT_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.550 296.000 138.830 300.000 ;
    END
  END DAT_O[31]
  PIN DAT_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 653.750 296.000 654.030 300.000 ;
    END
  END DAT_O[3]
  PIN DAT_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 663.410 296.000 663.690 300.000 ;
    END
  END DAT_O[4]
  PIN DAT_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 608.670 296.000 608.950 300.000 ;
    END
  END DAT_O[5]
  PIN DAT_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 631.210 296.000 631.490 300.000 ;
    END
  END DAT_O[6]
  PIN DAT_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 634.430 296.000 634.710 300.000 ;
    END
  END DAT_O[7]
  PIN DAT_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 476.650 296.000 476.930 300.000 ;
    END
  END DAT_O[8]
  PIN DAT_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 154.650 296.000 154.930 300.000 ;
    END
  END DAT_O[9]
  PIN SEL_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 296.000 109.850 300.000 ;
    END
  END SEL_O[0]
  PIN SEL_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 135.330 296.000 135.610 300.000 ;
    END
  END SEL_O[1]
  PIN SEL_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 199.730 296.000 200.010 300.000 ;
    END
  END SEL_O[2]
  PIN SEL_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 238.370 296.000 238.650 300.000 ;
    END
  END SEL_O[3]
  PIN STB_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.110 296.000 132.390 300.000 ;
    END
  END STB_O
  PIN WE_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 637.650 296.000 637.930 300.000 ;
    END
  END WE_O
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END clk
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 248.030 296.000 248.310 300.000 ;
    END
  END en
  PIN gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END gpio_in[0]
  PIN gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END gpio_in[10]
  PIN gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END gpio_in[11]
  PIN gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END gpio_in[12]
  PIN gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END gpio_in[13]
  PIN gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END gpio_in[14]
  PIN gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END gpio_in[15]
  PIN gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END gpio_in[16]
  PIN gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END gpio_in[17]
  PIN gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END gpio_in[18]
  PIN gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END gpio_in[19]
  PIN gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END gpio_in[1]
  PIN gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END gpio_in[20]
  PIN gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END gpio_in[21]
  PIN gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END gpio_in[22]
  PIN gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END gpio_in[23]
  PIN gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END gpio_in[24]
  PIN gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END gpio_in[25]
  PIN gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 157.870 296.000 158.150 300.000 ;
    END
  END gpio_in[26]
  PIN gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 215.830 296.000 216.110 300.000 ;
    END
  END gpio_in[27]
  PIN gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END gpio_in[28]
  PIN gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END gpio_in[29]
  PIN gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END gpio_in[2]
  PIN gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END gpio_in[30]
  PIN gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END gpio_in[31]
  PIN gpio_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END gpio_in[32]
  PIN gpio_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END gpio_in[33]
  PIN gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END gpio_in[3]
  PIN gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END gpio_in[4]
  PIN gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END gpio_in[5]
  PIN gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END gpio_in[6]
  PIN gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 444.450 296.000 444.730 300.000 ;
    END
  END gpio_in[7]
  PIN gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END gpio_in[8]
  PIN gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END gpio_in[9]
  PIN gpio_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 447.670 296.000 447.950 300.000 ;
    END
  END gpio_oeb[0]
  PIN gpio_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 296.000 129.170 300.000 ;
    END
  END gpio_oeb[10]
  PIN gpio_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 186.850 296.000 187.130 300.000 ;
    END
  END gpio_oeb[11]
  PIN gpio_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 241.590 296.000 241.870 300.000 ;
    END
  END gpio_oeb[12]
  PIN gpio_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 505.630 296.000 505.910 300.000 ;
    END
  END gpio_oeb[13]
  PIN gpio_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 528.170 296.000 528.450 300.000 ;
    END
  END gpio_oeb[14]
  PIN gpio_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 711.710 296.000 711.990 300.000 ;
    END
  END gpio_oeb[15]
  PIN gpio_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 656.970 296.000 657.250 300.000 ;
    END
  END gpio_oeb[16]
  PIN gpio_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 589.350 296.000 589.630 300.000 ;
    END
  END gpio_oeb[17]
  PIN gpio_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 708.490 296.000 708.770 300.000 ;
    END
  END gpio_oeb[18]
  PIN gpio_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 367.170 296.000 367.450 300.000 ;
    END
  END gpio_oeb[19]
  PIN gpio_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 363.950 296.000 364.230 300.000 ;
    END
  END gpio_oeb[1]
  PIN gpio_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 702.050 296.000 702.330 300.000 ;
    END
  END gpio_oeb[20]
  PIN gpio_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 721.370 296.000 721.650 300.000 ;
    END
  END gpio_oeb[21]
  PIN gpio_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 550.710 296.000 550.990 300.000 ;
    END
  END gpio_oeb[22]
  PIN gpio_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 296.000 125.950 300.000 ;
    END
  END gpio_oeb[23]
  PIN gpio_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 231.930 296.000 232.210 300.000 ;
    END
  END gpio_oeb[24]
  PIN gpio_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 296.000 106.630 300.000 ;
    END
  END gpio_oeb[25]
  PIN gpio_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 418.690 296.000 418.970 300.000 ;
    END
  END gpio_oeb[26]
  PIN gpio_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 225.490 296.000 225.770 300.000 ;
    END
  END gpio_oeb[27]
  PIN gpio_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 296.000 206.450 300.000 ;
    END
  END gpio_oeb[28]
  PIN gpio_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 164.310 296.000 164.590 300.000 ;
    END
  END gpio_oeb[29]
  PIN gpio_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 731.030 296.000 731.310 300.000 ;
    END
  END gpio_oeb[2]
  PIN gpio_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 170.750 296.000 171.030 300.000 ;
    END
  END gpio_oeb[30]
  PIN gpio_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 219.050 296.000 219.330 300.000 ;
    END
  END gpio_oeb[31]
  PIN gpio_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END gpio_oeb[32]
  PIN gpio_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END gpio_oeb[33]
  PIN gpio_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 647.310 296.000 647.590 300.000 ;
    END
  END gpio_oeb[3]
  PIN gpio_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 676.290 296.000 676.570 300.000 ;
    END
  END gpio_oeb[4]
  PIN gpio_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 724.590 296.000 724.870 300.000 ;
    END
  END gpio_oeb[5]
  PIN gpio_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 624.770 296.000 625.050 300.000 ;
    END
  END gpio_oeb[6]
  PIN gpio_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 650.530 296.000 650.810 300.000 ;
    END
  END gpio_oeb[7]
  PIN gpio_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 486.310 296.000 486.590 300.000 ;
    END
  END gpio_oeb[8]
  PIN gpio_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 296.000 122.730 300.000 ;
    END
  END gpio_oeb[9]
  PIN gpio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 392.930 296.000 393.210 300.000 ;
    END
  END gpio_out[0]
  PIN gpio_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 235.150 296.000 235.430 300.000 ;
    END
  END gpio_out[10]
  PIN gpio_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 193.290 296.000 193.570 300.000 ;
    END
  END gpio_out[11]
  PIN gpio_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 296.000 103.410 300.000 ;
    END
  END gpio_out[12]
  PIN gpio_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 508.850 296.000 509.130 300.000 ;
    END
  END gpio_out[13]
  PIN gpio_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 531.390 296.000 531.670 300.000 ;
    END
  END gpio_out[14]
  PIN gpio_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 714.930 296.000 715.210 300.000 ;
    END
  END gpio_out[15]
  PIN gpio_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 660.190 296.000 660.470 300.000 ;
    END
  END gpio_out[16]
  PIN gpio_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 586.130 296.000 586.410 300.000 ;
    END
  END gpio_out[17]
  PIN gpio_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 705.270 296.000 705.550 300.000 ;
    END
  END gpio_out[18]
  PIN gpio_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 370.390 296.000 370.670 300.000 ;
    END
  END gpio_out[19]
  PIN gpio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 360.730 296.000 361.010 300.000 ;
    END
  END gpio_out[1]
  PIN gpio_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 698.830 296.000 699.110 300.000 ;
    END
  END gpio_out[20]
  PIN gpio_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 718.150 296.000 718.430 300.000 ;
    END
  END gpio_out[21]
  PIN gpio_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 547.490 296.000 547.770 300.000 ;
    END
  END gpio_out[22]
  PIN gpio_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 177.190 296.000 177.470 300.000 ;
    END
  END gpio_out[23]
  PIN gpio_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 228.710 296.000 228.990 300.000 ;
    END
  END gpio_out[24]
  PIN gpio_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 202.950 296.000 203.230 300.000 ;
    END
  END gpio_out[25]
  PIN gpio_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 415.470 296.000 415.750 300.000 ;
    END
  END gpio_out[26]
  PIN gpio_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 209.390 296.000 209.670 300.000 ;
    END
  END gpio_out[27]
  PIN gpio_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 296.000 119.510 300.000 ;
    END
  END gpio_out[28]
  PIN gpio_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 296.000 100.190 300.000 ;
    END
  END gpio_out[29]
  PIN gpio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 734.250 296.000 734.530 300.000 ;
    END
  END gpio_out[2]
  PIN gpio_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 173.970 296.000 174.250 300.000 ;
    END
  END gpio_out[30]
  PIN gpio_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 296.000 93.750 300.000 ;
    END
  END gpio_out[31]
  PIN gpio_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END gpio_out[32]
  PIN gpio_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END gpio_out[33]
  PIN gpio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 644.090 296.000 644.370 300.000 ;
    END
  END gpio_out[3]
  PIN gpio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 673.070 296.000 673.350 300.000 ;
    END
  END gpio_out[4]
  PIN gpio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 727.810 296.000 728.090 300.000 ;
    END
  END gpio_out[5]
  PIN gpio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 621.550 296.000 621.830 300.000 ;
    END
  END gpio_out[6]
  PIN gpio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 640.870 296.000 641.150 300.000 ;
    END
  END gpio_out[7]
  PIN gpio_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 483.090 296.000 483.370 300.000 ;
    END
  END gpio_out[8]
  PIN gpio_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 161.090 296.000 161.370 300.000 ;
    END
  END gpio_out[9]
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 896.000 17.040 900.000 17.640 ;
    END
  END nrst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 10.640 793.940 288.560 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 894.430 288.405 ;
      LAYER li1 ;
        RECT 5.520 10.795 894.240 288.405 ;
      LAYER met1 ;
        RECT 5.520 6.500 894.240 291.000 ;
      LAYER met2 ;
        RECT 6.530 295.720 89.970 296.210 ;
        RECT 90.810 295.720 93.190 296.210 ;
        RECT 94.030 295.720 96.410 296.210 ;
        RECT 97.250 295.720 99.630 296.210 ;
        RECT 100.470 295.720 102.850 296.210 ;
        RECT 103.690 295.720 106.070 296.210 ;
        RECT 106.910 295.720 109.290 296.210 ;
        RECT 110.130 295.720 112.510 296.210 ;
        RECT 113.350 295.720 115.730 296.210 ;
        RECT 116.570 295.720 118.950 296.210 ;
        RECT 119.790 295.720 122.170 296.210 ;
        RECT 123.010 295.720 125.390 296.210 ;
        RECT 126.230 295.720 128.610 296.210 ;
        RECT 129.450 295.720 131.830 296.210 ;
        RECT 132.670 295.720 135.050 296.210 ;
        RECT 135.890 295.720 138.270 296.210 ;
        RECT 139.110 295.720 141.490 296.210 ;
        RECT 142.330 295.720 144.710 296.210 ;
        RECT 145.550 295.720 147.930 296.210 ;
        RECT 148.770 295.720 151.150 296.210 ;
        RECT 151.990 295.720 154.370 296.210 ;
        RECT 155.210 295.720 157.590 296.210 ;
        RECT 158.430 295.720 160.810 296.210 ;
        RECT 161.650 295.720 164.030 296.210 ;
        RECT 164.870 295.720 167.250 296.210 ;
        RECT 168.090 295.720 170.470 296.210 ;
        RECT 171.310 295.720 173.690 296.210 ;
        RECT 174.530 295.720 176.910 296.210 ;
        RECT 177.750 295.720 180.130 296.210 ;
        RECT 180.970 295.720 183.350 296.210 ;
        RECT 184.190 295.720 186.570 296.210 ;
        RECT 187.410 295.720 189.790 296.210 ;
        RECT 190.630 295.720 193.010 296.210 ;
        RECT 193.850 295.720 196.230 296.210 ;
        RECT 197.070 295.720 199.450 296.210 ;
        RECT 200.290 295.720 202.670 296.210 ;
        RECT 203.510 295.720 205.890 296.210 ;
        RECT 206.730 295.720 209.110 296.210 ;
        RECT 209.950 295.720 212.330 296.210 ;
        RECT 213.170 295.720 215.550 296.210 ;
        RECT 216.390 295.720 218.770 296.210 ;
        RECT 219.610 295.720 221.990 296.210 ;
        RECT 222.830 295.720 225.210 296.210 ;
        RECT 226.050 295.720 228.430 296.210 ;
        RECT 229.270 295.720 231.650 296.210 ;
        RECT 232.490 295.720 234.870 296.210 ;
        RECT 235.710 295.720 238.090 296.210 ;
        RECT 238.930 295.720 241.310 296.210 ;
        RECT 242.150 295.720 244.530 296.210 ;
        RECT 245.370 295.720 247.750 296.210 ;
        RECT 248.590 295.720 250.970 296.210 ;
        RECT 251.810 295.720 254.190 296.210 ;
        RECT 255.030 295.720 357.230 296.210 ;
        RECT 358.070 295.720 360.450 296.210 ;
        RECT 361.290 295.720 363.670 296.210 ;
        RECT 364.510 295.720 366.890 296.210 ;
        RECT 367.730 295.720 370.110 296.210 ;
        RECT 370.950 295.720 373.330 296.210 ;
        RECT 374.170 295.720 382.990 296.210 ;
        RECT 383.830 295.720 389.430 296.210 ;
        RECT 390.270 295.720 392.650 296.210 ;
        RECT 393.490 295.720 395.870 296.210 ;
        RECT 396.710 295.720 399.090 296.210 ;
        RECT 399.930 295.720 405.530 296.210 ;
        RECT 406.370 295.720 415.190 296.210 ;
        RECT 416.030 295.720 418.410 296.210 ;
        RECT 419.250 295.720 421.630 296.210 ;
        RECT 422.470 295.720 424.850 296.210 ;
        RECT 425.690 295.720 431.290 296.210 ;
        RECT 432.130 295.720 440.950 296.210 ;
        RECT 441.790 295.720 444.170 296.210 ;
        RECT 445.010 295.720 447.390 296.210 ;
        RECT 448.230 295.720 450.610 296.210 ;
        RECT 451.450 295.720 453.830 296.210 ;
        RECT 454.670 295.720 457.050 296.210 ;
        RECT 457.890 295.720 473.150 296.210 ;
        RECT 473.990 295.720 476.370 296.210 ;
        RECT 477.210 295.720 479.590 296.210 ;
        RECT 480.430 295.720 482.810 296.210 ;
        RECT 483.650 295.720 486.030 296.210 ;
        RECT 486.870 295.720 489.250 296.210 ;
        RECT 490.090 295.720 502.130 296.210 ;
        RECT 502.970 295.720 505.350 296.210 ;
        RECT 506.190 295.720 508.570 296.210 ;
        RECT 509.410 295.720 511.790 296.210 ;
        RECT 512.630 295.720 524.670 296.210 ;
        RECT 525.510 295.720 527.890 296.210 ;
        RECT 528.730 295.720 531.110 296.210 ;
        RECT 531.950 295.720 534.330 296.210 ;
        RECT 535.170 295.720 537.550 296.210 ;
        RECT 538.390 295.720 540.770 296.210 ;
        RECT 541.610 295.720 547.210 296.210 ;
        RECT 548.050 295.720 550.430 296.210 ;
        RECT 551.270 295.720 556.870 296.210 ;
        RECT 557.710 295.720 560.090 296.210 ;
        RECT 560.930 295.720 563.310 296.210 ;
        RECT 564.150 295.720 572.970 296.210 ;
        RECT 573.810 295.720 576.190 296.210 ;
        RECT 577.030 295.720 579.410 296.210 ;
        RECT 580.250 295.720 585.850 296.210 ;
        RECT 586.690 295.720 589.070 296.210 ;
        RECT 589.910 295.720 592.290 296.210 ;
        RECT 593.130 295.720 595.510 296.210 ;
        RECT 596.350 295.720 608.390 296.210 ;
        RECT 609.230 295.720 611.610 296.210 ;
        RECT 612.450 295.720 614.830 296.210 ;
        RECT 615.670 295.720 618.050 296.210 ;
        RECT 618.890 295.720 621.270 296.210 ;
        RECT 622.110 295.720 624.490 296.210 ;
        RECT 625.330 295.720 630.930 296.210 ;
        RECT 631.770 295.720 634.150 296.210 ;
        RECT 634.990 295.720 637.370 296.210 ;
        RECT 638.210 295.720 640.590 296.210 ;
        RECT 641.430 295.720 643.810 296.210 ;
        RECT 644.650 295.720 647.030 296.210 ;
        RECT 647.870 295.720 650.250 296.210 ;
        RECT 651.090 295.720 653.470 296.210 ;
        RECT 654.310 295.720 656.690 296.210 ;
        RECT 657.530 295.720 659.910 296.210 ;
        RECT 660.750 295.720 663.130 296.210 ;
        RECT 663.970 295.720 666.350 296.210 ;
        RECT 667.190 295.720 669.570 296.210 ;
        RECT 670.410 295.720 672.790 296.210 ;
        RECT 673.630 295.720 676.010 296.210 ;
        RECT 676.850 295.720 685.670 296.210 ;
        RECT 686.510 295.720 688.890 296.210 ;
        RECT 689.730 295.720 692.110 296.210 ;
        RECT 692.950 295.720 695.330 296.210 ;
        RECT 696.170 295.720 698.550 296.210 ;
        RECT 699.390 295.720 701.770 296.210 ;
        RECT 702.610 295.720 704.990 296.210 ;
        RECT 705.830 295.720 708.210 296.210 ;
        RECT 709.050 295.720 711.430 296.210 ;
        RECT 712.270 295.720 714.650 296.210 ;
        RECT 715.490 295.720 717.870 296.210 ;
        RECT 718.710 295.720 721.090 296.210 ;
        RECT 721.930 295.720 724.310 296.210 ;
        RECT 725.150 295.720 727.530 296.210 ;
        RECT 728.370 295.720 730.750 296.210 ;
        RECT 731.590 295.720 733.970 296.210 ;
        RECT 734.810 295.720 892.770 296.210 ;
        RECT 6.530 4.280 892.770 295.720 ;
        RECT 6.530 0.155 25.570 4.280 ;
        RECT 26.410 0.155 247.750 4.280 ;
        RECT 248.590 0.155 250.970 4.280 ;
        RECT 251.810 0.155 254.190 4.280 ;
        RECT 255.030 0.155 257.410 4.280 ;
        RECT 258.250 0.155 260.630 4.280 ;
        RECT 261.470 0.155 263.850 4.280 ;
        RECT 264.690 0.155 267.070 4.280 ;
        RECT 267.910 0.155 270.290 4.280 ;
        RECT 271.130 0.155 273.510 4.280 ;
        RECT 274.350 0.155 276.730 4.280 ;
        RECT 277.570 0.155 279.950 4.280 ;
        RECT 280.790 0.155 283.170 4.280 ;
        RECT 284.010 0.155 286.390 4.280 ;
        RECT 287.230 0.155 289.610 4.280 ;
        RECT 290.450 0.155 292.830 4.280 ;
        RECT 293.670 0.155 296.050 4.280 ;
        RECT 296.890 0.155 299.270 4.280 ;
        RECT 300.110 0.155 302.490 4.280 ;
        RECT 303.330 0.155 305.710 4.280 ;
        RECT 306.550 0.155 308.930 4.280 ;
        RECT 309.770 0.155 312.150 4.280 ;
        RECT 312.990 0.155 315.370 4.280 ;
        RECT 316.210 0.155 318.590 4.280 ;
        RECT 319.430 0.155 321.810 4.280 ;
        RECT 322.650 0.155 325.030 4.280 ;
        RECT 325.870 0.155 328.250 4.280 ;
        RECT 329.090 0.155 331.470 4.280 ;
        RECT 332.310 0.155 334.690 4.280 ;
        RECT 335.530 0.155 337.910 4.280 ;
        RECT 338.750 0.155 341.130 4.280 ;
        RECT 341.970 0.155 344.350 4.280 ;
        RECT 345.190 0.155 347.570 4.280 ;
        RECT 348.410 0.155 350.790 4.280 ;
        RECT 351.630 0.155 354.010 4.280 ;
        RECT 354.850 0.155 357.230 4.280 ;
        RECT 358.070 0.155 360.450 4.280 ;
        RECT 361.290 0.155 363.670 4.280 ;
        RECT 364.510 0.155 366.890 4.280 ;
        RECT 367.730 0.155 370.110 4.280 ;
        RECT 370.950 0.155 373.330 4.280 ;
        RECT 374.170 0.155 376.550 4.280 ;
        RECT 377.390 0.155 379.770 4.280 ;
        RECT 380.610 0.155 382.990 4.280 ;
        RECT 383.830 0.155 386.210 4.280 ;
        RECT 387.050 0.155 389.430 4.280 ;
        RECT 390.270 0.155 392.650 4.280 ;
        RECT 393.490 0.155 395.870 4.280 ;
        RECT 396.710 0.155 399.090 4.280 ;
        RECT 399.930 0.155 402.310 4.280 ;
        RECT 403.150 0.155 405.530 4.280 ;
        RECT 406.370 0.155 408.750 4.280 ;
        RECT 409.590 0.155 411.970 4.280 ;
        RECT 412.810 0.155 415.190 4.280 ;
        RECT 416.030 0.155 418.410 4.280 ;
        RECT 419.250 0.155 424.850 4.280 ;
        RECT 425.690 0.155 431.290 4.280 ;
        RECT 432.130 0.155 434.510 4.280 ;
        RECT 435.350 0.155 437.730 4.280 ;
        RECT 438.570 0.155 440.950 4.280 ;
        RECT 441.790 0.155 450.610 4.280 ;
        RECT 451.450 0.155 453.830 4.280 ;
        RECT 454.670 0.155 892.770 4.280 ;
      LAYER met3 ;
        RECT 4.000 266.240 896.000 290.185 ;
        RECT 4.400 264.840 896.000 266.240 ;
        RECT 4.000 262.840 896.000 264.840 ;
        RECT 4.400 261.440 896.000 262.840 ;
        RECT 4.000 259.440 896.000 261.440 ;
        RECT 4.400 258.040 896.000 259.440 ;
        RECT 4.000 256.040 896.000 258.040 ;
        RECT 4.400 254.640 896.000 256.040 ;
        RECT 4.000 18.040 896.000 254.640 ;
        RECT 4.000 16.640 895.600 18.040 ;
        RECT 4.000 0.175 896.000 16.640 ;
      LAYER met4 ;
        RECT 35.255 288.960 881.065 290.185 ;
        RECT 35.255 10.240 174.240 288.960 ;
        RECT 176.640 10.240 177.540 288.960 ;
        RECT 179.940 10.240 327.840 288.960 ;
        RECT 330.240 10.240 331.140 288.960 ;
        RECT 333.540 10.240 481.440 288.960 ;
        RECT 483.840 10.240 484.740 288.960 ;
        RECT 487.140 10.240 635.040 288.960 ;
        RECT 637.440 10.240 638.340 288.960 ;
        RECT 640.740 10.240 788.640 288.960 ;
        RECT 791.040 10.240 791.940 288.960 ;
        RECT 794.340 10.240 881.065 288.960 ;
        RECT 35.255 0.175 881.065 10.240 ;
  END
END team_03
END LIBRARY

